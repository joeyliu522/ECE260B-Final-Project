##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 15:55:39 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1260.0000 BY 1720.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1000.0500 0.0000 1000.1500 0.5200 ;
    END
  END clk
  PIN sum_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 860.1500 0.5200 860.2500 ;
    END
  END sum_in[23]
  PIN sum_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 865.1500 0.5200 865.2500 ;
    END
  END sum_in[22]
  PIN sum_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 870.1500 0.5200 870.2500 ;
    END
  END sum_in[21]
  PIN sum_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 875.1500 0.5200 875.2500 ;
    END
  END sum_in[20]
  PIN sum_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 880.1500 0.5200 880.2500 ;
    END
  END sum_in[19]
  PIN sum_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 885.1500 0.5200 885.2500 ;
    END
  END sum_in[18]
  PIN sum_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 890.1500 0.5200 890.2500 ;
    END
  END sum_in[17]
  PIN sum_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 895.1500 0.5200 895.2500 ;
    END
  END sum_in[16]
  PIN sum_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 900.1500 0.5200 900.2500 ;
    END
  END sum_in[15]
  PIN sum_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 905.1500 0.5200 905.2500 ;
    END
  END sum_in[14]
  PIN sum_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 910.1500 0.5200 910.2500 ;
    END
  END sum_in[13]
  PIN sum_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 915.1500 0.5200 915.2500 ;
    END
  END sum_in[12]
  PIN sum_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 920.1500 0.5200 920.2500 ;
    END
  END sum_in[11]
  PIN sum_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 925.1500 0.5200 925.2500 ;
    END
  END sum_in[10]
  PIN sum_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 930.1500 0.5200 930.2500 ;
    END
  END sum_in[9]
  PIN sum_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 935.1500 0.5200 935.2500 ;
    END
  END sum_in[8]
  PIN sum_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 940.1500 0.5200 940.2500 ;
    END
  END sum_in[7]
  PIN sum_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 945.1500 0.5200 945.2500 ;
    END
  END sum_in[6]
  PIN sum_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 950.1500 0.5200 950.2500 ;
    END
  END sum_in[5]
  PIN sum_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 955.1500 0.5200 955.2500 ;
    END
  END sum_in[4]
  PIN sum_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 960.1500 0.5200 960.2500 ;
    END
  END sum_in[3]
  PIN sum_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 965.1500 0.5200 965.2500 ;
    END
  END sum_in[2]
  PIN sum_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 970.1500 0.5200 970.2500 ;
    END
  END sum_in[1]
  PIN sum_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 975.1500 0.5200 975.2500 ;
    END
  END sum_in[0]
  PIN fifo_ext_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 980.1500 0.5200 980.2500 ;
    END
  END fifo_ext_rd
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 740.1500 0.5200 740.2500 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 745.1500 0.5200 745.2500 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 750.1500 0.5200 750.2500 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 755.1500 0.5200 755.2500 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 760.1500 0.5200 760.2500 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 765.1500 0.5200 765.2500 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 770.1500 0.5200 770.2500 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 775.1500 0.5200 775.2500 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 780.1500 0.5200 780.2500 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 785.1500 0.5200 785.2500 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 790.1500 0.5200 790.2500 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 795.1500 0.5200 795.2500 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 800.1500 0.5200 800.2500 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 805.1500 0.5200 805.2500 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 810.1500 0.5200 810.2500 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 815.1500 0.5200 815.2500 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 820.1500 0.5200 820.2500 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 825.1500 0.5200 825.2500 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 830.1500 0.5200 830.2500 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 835.1500 0.5200 835.2500 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 840.1500 0.5200 840.2500 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 845.1500 0.5200 845.2500 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 850.1500 0.5200 850.2500 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 855.1500 0.5200 855.2500 ;
    END
  END sum_out[0]
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.0500 0.0000 260.1500 0.5200 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.0500 0.0000 265.1500 0.5200 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.0500 0.0000 270.1500 0.5200 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.0500 0.0000 275.1500 0.5200 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.0500 0.0000 280.1500 0.5200 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.0500 0.0000 285.1500 0.5200 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.0500 0.0000 290.1500 0.5200 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.0500 0.0000 295.1500 0.5200 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.0500 0.0000 300.1500 0.5200 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.0500 0.0000 305.1500 0.5200 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.0500 0.0000 310.1500 0.5200 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.0500 0.0000 315.1500 0.5200 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.0500 0.0000 320.1500 0.5200 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.0500 0.0000 325.1500 0.5200 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.0500 0.0000 330.1500 0.5200 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.0500 0.0000 335.1500 0.5200 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.0500 0.0000 340.1500 0.5200 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.0500 0.0000 345.1500 0.5200 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.0500 0.0000 350.1500 0.5200 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.0500 0.0000 355.1500 0.5200 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.0500 0.0000 360.1500 0.5200 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.0500 0.0000 365.1500 0.5200 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.0500 0.0000 370.1500 0.5200 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.0500 0.0000 375.1500 0.5200 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.0500 0.0000 380.1500 0.5200 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.0500 0.0000 385.1500 0.5200 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.0500 0.0000 390.1500 0.5200 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.0500 0.0000 395.1500 0.5200 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.0500 0.0000 400.1500 0.5200 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.0500 0.0000 405.1500 0.5200 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.0500 0.0000 410.1500 0.5200 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.0500 0.0000 415.1500 0.5200 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.0500 0.0000 420.1500 0.5200 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.0500 0.0000 425.1500 0.5200 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.0500 0.0000 430.1500 0.5200 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.0500 0.0000 435.1500 0.5200 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.0500 0.0000 440.1500 0.5200 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.0500 0.0000 445.1500 0.5200 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.0500 0.0000 450.1500 0.5200 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.0500 0.0000 455.1500 0.5200 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.0500 0.0000 460.1500 0.5200 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 465.0500 0.0000 465.1500 0.5200 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.0500 0.0000 470.1500 0.5200 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.0500 0.0000 475.1500 0.5200 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 480.0500 0.0000 480.1500 0.5200 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.0500 0.0000 485.1500 0.5200 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 490.0500 0.0000 490.1500 0.5200 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.0500 0.0000 495.1500 0.5200 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.0500 0.0000 500.1500 0.5200 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 505.0500 0.0000 505.1500 0.5200 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.0500 0.0000 510.1500 0.5200 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.0500 0.0000 515.1500 0.5200 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 520.0500 0.0000 520.1500 0.5200 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.0500 0.0000 525.1500 0.5200 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 530.0500 0.0000 530.1500 0.5200 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.0500 0.0000 535.1500 0.5200 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 540.0500 0.0000 540.1500 0.5200 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 545.0500 0.0000 545.1500 0.5200 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 550.0500 0.0000 550.1500 0.5200 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.0500 0.0000 555.1500 0.5200 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 560.0500 0.0000 560.1500 0.5200 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.0500 0.0000 565.1500 0.5200 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 570.0500 0.0000 570.1500 0.5200 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.0500 0.0000 575.1500 0.5200 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 580.0500 0.0000 580.1500 0.5200 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 585.0500 0.0000 585.1500 0.5200 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 590.0500 0.0000 590.1500 0.5200 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.0500 0.0000 595.1500 0.5200 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 600.0500 0.0000 600.1500 0.5200 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 605.0500 0.0000 605.1500 0.5200 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 610.0500 0.0000 610.1500 0.5200 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.0500 0.0000 615.1500 0.5200 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 620.0500 0.0000 620.1500 0.5200 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 625.0500 0.0000 625.1500 0.5200 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 630.0500 0.0000 630.1500 0.5200 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.0500 0.0000 635.1500 0.5200 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 640.0500 0.0000 640.1500 0.5200 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 645.0500 0.0000 645.1500 0.5200 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 650.0500 0.0000 650.1500 0.5200 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.0500 0.0000 655.1500 0.5200 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 660.0500 0.0000 660.1500 0.5200 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.0500 0.0000 665.1500 0.5200 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 670.0500 0.0000 670.1500 0.5200 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.0500 0.0000 675.1500 0.5200 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 680.0500 0.0000 680.1500 0.5200 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 685.0500 0.0000 685.1500 0.5200 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690.0500 0.0000 690.1500 0.5200 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 695.0500 0.0000 695.1500 0.5200 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 700.0500 0.0000 700.1500 0.5200 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 705.0500 0.0000 705.1500 0.5200 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 710.0500 0.0000 710.1500 0.5200 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 715.0500 0.0000 715.1500 0.5200 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 720.0500 0.0000 720.1500 0.5200 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 725.0500 0.0000 725.1500 0.5200 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 730.0500 0.0000 730.1500 0.5200 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 735.0500 0.0000 735.1500 0.5200 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 740.0500 0.0000 740.1500 0.5200 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 745.0500 0.0000 745.1500 0.5200 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 750.0500 0.0000 750.1500 0.5200 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 755.0500 0.0000 755.1500 0.5200 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 760.0500 0.0000 760.1500 0.5200 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 765.0500 0.0000 765.1500 0.5200 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 770.0500 0.0000 770.1500 0.5200 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 775.0500 0.0000 775.1500 0.5200 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 780.0500 0.0000 780.1500 0.5200 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 785.0500 0.0000 785.1500 0.5200 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 790.0500 0.0000 790.1500 0.5200 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 795.0500 0.0000 795.1500 0.5200 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 800.0500 0.0000 800.1500 0.5200 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 805.0500 0.0000 805.1500 0.5200 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 810.0500 0.0000 810.1500 0.5200 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 815.0500 0.0000 815.1500 0.5200 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 820.0500 0.0000 820.1500 0.5200 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 825.0500 0.0000 825.1500 0.5200 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 830.0500 0.0000 830.1500 0.5200 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 835.0500 0.0000 835.1500 0.5200 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 840.0500 0.0000 840.1500 0.5200 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 845.0500 0.0000 845.1500 0.5200 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 850.0500 0.0000 850.1500 0.5200 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 855.0500 0.0000 855.1500 0.5200 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 860.0500 0.0000 860.1500 0.5200 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 865.0500 0.0000 865.1500 0.5200 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 870.0500 0.0000 870.1500 0.5200 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 875.0500 0.0000 875.1500 0.5200 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 880.0500 0.0000 880.1500 0.5200 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 885.0500 0.0000 885.1500 0.5200 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 890.0500 0.0000 890.1500 0.5200 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 895.0500 0.0000 895.1500 0.5200 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1027.2500 1719.4800 1027.3500 1720.0000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1022.2500 1719.4800 1022.3500 1720.0000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1017.2500 1719.4800 1017.3500 1720.0000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1012.2500 1719.4800 1012.3500 1720.0000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1007.2500 1719.4800 1007.3500 1720.0000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1002.2500 1719.4800 1002.3500 1720.0000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 997.2500 1719.4800 997.3500 1720.0000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 992.2500 1719.4800 992.3500 1720.0000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 987.2500 1719.4800 987.3500 1720.0000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 982.2500 1719.4800 982.3500 1720.0000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 977.2500 1719.4800 977.3500 1720.0000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 972.2500 1719.4800 972.3500 1720.0000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 967.2500 1719.4800 967.3500 1720.0000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 962.2500 1719.4800 962.3500 1720.0000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 957.2500 1719.4800 957.3500 1720.0000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 952.2500 1719.4800 952.3500 1720.0000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 947.2500 1719.4800 947.3500 1720.0000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 942.2500 1719.4800 942.3500 1720.0000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 937.2500 1719.4800 937.3500 1720.0000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 932.2500 1719.4800 932.3500 1720.0000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 927.2500 1719.4800 927.3500 1720.0000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 922.2500 1719.4800 922.3500 1720.0000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 917.2500 1719.4800 917.3500 1720.0000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 912.2500 1719.4800 912.3500 1720.0000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 907.2500 1719.4800 907.3500 1720.0000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 902.2500 1719.4800 902.3500 1720.0000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 897.2500 1719.4800 897.3500 1720.0000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 892.2500 1719.4800 892.3500 1720.0000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 887.2500 1719.4800 887.3500 1720.0000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 882.2500 1719.4800 882.3500 1720.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 877.2500 1719.4800 877.3500 1720.0000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 872.2500 1719.4800 872.3500 1720.0000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 867.2500 1719.4800 867.3500 1720.0000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 862.2500 1719.4800 862.3500 1720.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 857.2500 1719.4800 857.3500 1720.0000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 852.2500 1719.4800 852.3500 1720.0000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 847.2500 1719.4800 847.3500 1720.0000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 842.2500 1719.4800 842.3500 1720.0000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 837.2500 1719.4800 837.3500 1720.0000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 832.2500 1719.4800 832.3500 1720.0000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 827.2500 1719.4800 827.3500 1720.0000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 822.2500 1719.4800 822.3500 1720.0000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 817.2500 1719.4800 817.3500 1720.0000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 812.2500 1719.4800 812.3500 1720.0000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 807.2500 1719.4800 807.3500 1720.0000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 802.2500 1719.4800 802.3500 1720.0000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 797.2500 1719.4800 797.3500 1720.0000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 792.2500 1719.4800 792.3500 1720.0000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 787.2500 1719.4800 787.3500 1720.0000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 782.2500 1719.4800 782.3500 1720.0000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 777.2500 1719.4800 777.3500 1720.0000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 772.2500 1719.4800 772.3500 1720.0000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 767.2500 1719.4800 767.3500 1720.0000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 762.2500 1719.4800 762.3500 1720.0000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 757.2500 1719.4800 757.3500 1720.0000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 752.2500 1719.4800 752.3500 1720.0000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 747.2500 1719.4800 747.3500 1720.0000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 742.2500 1719.4800 742.3500 1720.0000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 737.2500 1719.4800 737.3500 1720.0000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 732.2500 1719.4800 732.3500 1720.0000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 727.2500 1719.4800 727.3500 1720.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 722.2500 1719.4800 722.3500 1720.0000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 717.2500 1719.4800 717.3500 1720.0000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 712.2500 1719.4800 712.3500 1720.0000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 707.2500 1719.4800 707.3500 1720.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 702.2500 1719.4800 702.3500 1720.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 697.2500 1719.4800 697.3500 1720.0000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 692.2500 1719.4800 692.3500 1720.0000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.2500 1719.4800 687.3500 1720.0000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 682.2500 1719.4800 682.3500 1720.0000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 677.2500 1719.4800 677.3500 1720.0000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 672.2500 1719.4800 672.3500 1720.0000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.2500 1719.4800 667.3500 1720.0000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 662.2500 1719.4800 662.3500 1720.0000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 657.2500 1719.4800 657.3500 1720.0000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 652.2500 1719.4800 652.3500 1720.0000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.2500 1719.4800 647.3500 1720.0000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 642.2500 1719.4800 642.3500 1720.0000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 637.2500 1719.4800 637.3500 1720.0000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 632.2500 1719.4800 632.3500 1720.0000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.2500 1719.4800 627.3500 1720.0000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 622.2500 1719.4800 622.3500 1720.0000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 617.2500 1719.4800 617.3500 1720.0000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 612.2500 1719.4800 612.3500 1720.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.2500 1719.4800 607.3500 1720.0000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 602.2500 1719.4800 602.3500 1720.0000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 597.2500 1719.4800 597.3500 1720.0000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 592.2500 1719.4800 592.3500 1720.0000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.2500 1719.4800 587.3500 1720.0000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 582.2500 1719.4800 582.3500 1720.0000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 577.2500 1719.4800 577.3500 1720.0000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.2500 1719.4800 572.3500 1720.0000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.2500 1719.4800 567.3500 1720.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 562.2500 1719.4800 562.3500 1720.0000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 557.2500 1719.4800 557.3500 1720.0000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 552.2500 1719.4800 552.3500 1720.0000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.2500 1719.4800 547.3500 1720.0000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 542.2500 1719.4800 542.3500 1720.0000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 537.2500 1719.4800 537.3500 1720.0000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 532.2500 1719.4800 532.3500 1720.0000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.2500 1719.4800 527.3500 1720.0000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 522.2500 1719.4800 522.3500 1720.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 517.2500 1719.4800 517.3500 1720.0000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 512.2500 1719.4800 512.3500 1720.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.2500 1719.4800 507.3500 1720.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 502.2500 1719.4800 502.3500 1720.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.2500 1719.4800 497.3500 1720.0000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.2500 1719.4800 492.3500 1720.0000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.2500 1719.4800 487.3500 1720.0000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 482.2500 1719.4800 482.3500 1720.0000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.2500 1719.4800 477.3500 1720.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 472.2500 1719.4800 472.3500 1720.0000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.2500 1719.4800 467.3500 1720.0000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 462.2500 1719.4800 462.3500 1720.0000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.2500 1719.4800 457.3500 1720.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.2500 1719.4800 452.3500 1720.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.2500 1719.4800 447.3500 1720.0000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.2500 1719.4800 442.3500 1720.0000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.2500 1719.4800 437.3500 1720.0000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.2500 1719.4800 432.3500 1720.0000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.2500 1719.4800 427.3500 1720.0000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.2500 1719.4800 422.3500 1720.0000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.2500 1719.4800 417.3500 1720.0000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.2500 1719.4800 412.3500 1720.0000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.2500 1719.4800 407.3500 1720.0000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.2500 1719.4800 402.3500 1720.0000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.2500 1719.4800 397.3500 1720.0000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.2500 1719.4800 392.3500 1720.0000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.2500 1719.4800 387.3500 1720.0000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.2500 1719.4800 382.3500 1720.0000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.2500 1719.4800 377.3500 1720.0000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.2500 1719.4800 372.3500 1720.0000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.2500 1719.4800 367.3500 1720.0000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.2500 1719.4800 362.3500 1720.0000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.2500 1719.4800 357.3500 1720.0000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.2500 1719.4800 352.3500 1720.0000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.2500 1719.4800 347.3500 1720.0000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.2500 1719.4800 342.3500 1720.0000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.2500 1719.4800 337.3500 1720.0000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.2500 1719.4800 332.3500 1720.0000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.2500 1719.4800 327.3500 1720.0000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.2500 1719.4800 322.3500 1720.0000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.2500 1719.4800 317.3500 1720.0000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.2500 1719.4800 312.3500 1720.0000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.2500 1719.4800 307.3500 1720.0000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.2500 1719.4800 302.3500 1720.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.2500 1719.4800 297.3500 1720.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.2500 1719.4800 292.3500 1720.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.2500 1719.4800 287.3500 1720.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.2500 1719.4800 282.3500 1720.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.2500 1719.4800 277.3500 1720.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.2500 1719.4800 272.3500 1720.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.2500 1719.4800 267.3500 1720.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.2500 1719.4800 262.3500 1720.0000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.2500 1719.4800 257.3500 1720.0000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.2500 1719.4800 252.3500 1720.0000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.2500 1719.4800 247.3500 1720.0000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.2500 1719.4800 242.3500 1720.0000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.2500 1719.4800 237.3500 1720.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.2500 1719.4800 232.3500 1720.0000 ;
    END
  END out[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 900.0500 0.0000 900.1500 0.5200 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 905.0500 0.0000 905.1500 0.5200 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 910.0500 0.0000 910.1500 0.5200 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 915.0500 0.0000 915.1500 0.5200 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 920.0500 0.0000 920.1500 0.5200 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 925.0500 0.0000 925.1500 0.5200 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 930.0500 0.0000 930.1500 0.5200 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 935.0500 0.0000 935.1500 0.5200 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 940.0500 0.0000 940.1500 0.5200 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 945.0500 0.0000 945.1500 0.5200 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 950.0500 0.0000 950.1500 0.5200 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 955.0500 0.0000 955.1500 0.5200 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 960.0500 0.0000 960.1500 0.5200 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 965.0500 0.0000 965.1500 0.5200 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 970.0500 0.0000 970.1500 0.5200 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 975.0500 0.0000 975.1500 0.5200 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 980.0500 0.0000 980.1500 0.5200 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 985.0500 0.0000 985.1500 0.5200 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 990.0500 0.0000 990.1500 0.5200 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 995.0500 0.0000 995.1500 0.5200 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
    LAYER M2 ;
      RECT 1027.4500 1719.3800 1260.0000 1720.0000 ;
      RECT 1022.4500 1719.3800 1027.1500 1720.0000 ;
      RECT 1017.4500 1719.3800 1022.1500 1720.0000 ;
      RECT 1012.4500 1719.3800 1017.1500 1720.0000 ;
      RECT 1007.4500 1719.3800 1012.1500 1720.0000 ;
      RECT 1002.4500 1719.3800 1007.1500 1720.0000 ;
      RECT 997.4500 1719.3800 1002.1500 1720.0000 ;
      RECT 992.4500 1719.3800 997.1500 1720.0000 ;
      RECT 987.4500 1719.3800 992.1500 1720.0000 ;
      RECT 982.4500 1719.3800 987.1500 1720.0000 ;
      RECT 977.4500 1719.3800 982.1500 1720.0000 ;
      RECT 972.4500 1719.3800 977.1500 1720.0000 ;
      RECT 967.4500 1719.3800 972.1500 1720.0000 ;
      RECT 962.4500 1719.3800 967.1500 1720.0000 ;
      RECT 957.4500 1719.3800 962.1500 1720.0000 ;
      RECT 952.4500 1719.3800 957.1500 1720.0000 ;
      RECT 947.4500 1719.3800 952.1500 1720.0000 ;
      RECT 942.4500 1719.3800 947.1500 1720.0000 ;
      RECT 937.4500 1719.3800 942.1500 1720.0000 ;
      RECT 932.4500 1719.3800 937.1500 1720.0000 ;
      RECT 927.4500 1719.3800 932.1500 1720.0000 ;
      RECT 922.4500 1719.3800 927.1500 1720.0000 ;
      RECT 917.4500 1719.3800 922.1500 1720.0000 ;
      RECT 912.4500 1719.3800 917.1500 1720.0000 ;
      RECT 907.4500 1719.3800 912.1500 1720.0000 ;
      RECT 902.4500 1719.3800 907.1500 1720.0000 ;
      RECT 897.4500 1719.3800 902.1500 1720.0000 ;
      RECT 892.4500 1719.3800 897.1500 1720.0000 ;
      RECT 887.4500 1719.3800 892.1500 1720.0000 ;
      RECT 882.4500 1719.3800 887.1500 1720.0000 ;
      RECT 877.4500 1719.3800 882.1500 1720.0000 ;
      RECT 872.4500 1719.3800 877.1500 1720.0000 ;
      RECT 867.4500 1719.3800 872.1500 1720.0000 ;
      RECT 862.4500 1719.3800 867.1500 1720.0000 ;
      RECT 857.4500 1719.3800 862.1500 1720.0000 ;
      RECT 852.4500 1719.3800 857.1500 1720.0000 ;
      RECT 847.4500 1719.3800 852.1500 1720.0000 ;
      RECT 842.4500 1719.3800 847.1500 1720.0000 ;
      RECT 837.4500 1719.3800 842.1500 1720.0000 ;
      RECT 832.4500 1719.3800 837.1500 1720.0000 ;
      RECT 827.4500 1719.3800 832.1500 1720.0000 ;
      RECT 822.4500 1719.3800 827.1500 1720.0000 ;
      RECT 817.4500 1719.3800 822.1500 1720.0000 ;
      RECT 812.4500 1719.3800 817.1500 1720.0000 ;
      RECT 807.4500 1719.3800 812.1500 1720.0000 ;
      RECT 802.4500 1719.3800 807.1500 1720.0000 ;
      RECT 797.4500 1719.3800 802.1500 1720.0000 ;
      RECT 792.4500 1719.3800 797.1500 1720.0000 ;
      RECT 787.4500 1719.3800 792.1500 1720.0000 ;
      RECT 782.4500 1719.3800 787.1500 1720.0000 ;
      RECT 777.4500 1719.3800 782.1500 1720.0000 ;
      RECT 772.4500 1719.3800 777.1500 1720.0000 ;
      RECT 767.4500 1719.3800 772.1500 1720.0000 ;
      RECT 762.4500 1719.3800 767.1500 1720.0000 ;
      RECT 757.4500 1719.3800 762.1500 1720.0000 ;
      RECT 752.4500 1719.3800 757.1500 1720.0000 ;
      RECT 747.4500 1719.3800 752.1500 1720.0000 ;
      RECT 742.4500 1719.3800 747.1500 1720.0000 ;
      RECT 737.4500 1719.3800 742.1500 1720.0000 ;
      RECT 732.4500 1719.3800 737.1500 1720.0000 ;
      RECT 727.4500 1719.3800 732.1500 1720.0000 ;
      RECT 722.4500 1719.3800 727.1500 1720.0000 ;
      RECT 717.4500 1719.3800 722.1500 1720.0000 ;
      RECT 712.4500 1719.3800 717.1500 1720.0000 ;
      RECT 707.4500 1719.3800 712.1500 1720.0000 ;
      RECT 702.4500 1719.3800 707.1500 1720.0000 ;
      RECT 697.4500 1719.3800 702.1500 1720.0000 ;
      RECT 692.4500 1719.3800 697.1500 1720.0000 ;
      RECT 687.4500 1719.3800 692.1500 1720.0000 ;
      RECT 682.4500 1719.3800 687.1500 1720.0000 ;
      RECT 677.4500 1719.3800 682.1500 1720.0000 ;
      RECT 672.4500 1719.3800 677.1500 1720.0000 ;
      RECT 667.4500 1719.3800 672.1500 1720.0000 ;
      RECT 662.4500 1719.3800 667.1500 1720.0000 ;
      RECT 657.4500 1719.3800 662.1500 1720.0000 ;
      RECT 652.4500 1719.3800 657.1500 1720.0000 ;
      RECT 647.4500 1719.3800 652.1500 1720.0000 ;
      RECT 642.4500 1719.3800 647.1500 1720.0000 ;
      RECT 637.4500 1719.3800 642.1500 1720.0000 ;
      RECT 632.4500 1719.3800 637.1500 1720.0000 ;
      RECT 627.4500 1719.3800 632.1500 1720.0000 ;
      RECT 622.4500 1719.3800 627.1500 1720.0000 ;
      RECT 617.4500 1719.3800 622.1500 1720.0000 ;
      RECT 612.4500 1719.3800 617.1500 1720.0000 ;
      RECT 607.4500 1719.3800 612.1500 1720.0000 ;
      RECT 602.4500 1719.3800 607.1500 1720.0000 ;
      RECT 597.4500 1719.3800 602.1500 1720.0000 ;
      RECT 592.4500 1719.3800 597.1500 1720.0000 ;
      RECT 587.4500 1719.3800 592.1500 1720.0000 ;
      RECT 582.4500 1719.3800 587.1500 1720.0000 ;
      RECT 577.4500 1719.3800 582.1500 1720.0000 ;
      RECT 572.4500 1719.3800 577.1500 1720.0000 ;
      RECT 567.4500 1719.3800 572.1500 1720.0000 ;
      RECT 562.4500 1719.3800 567.1500 1720.0000 ;
      RECT 557.4500 1719.3800 562.1500 1720.0000 ;
      RECT 552.4500 1719.3800 557.1500 1720.0000 ;
      RECT 547.4500 1719.3800 552.1500 1720.0000 ;
      RECT 542.4500 1719.3800 547.1500 1720.0000 ;
      RECT 537.4500 1719.3800 542.1500 1720.0000 ;
      RECT 532.4500 1719.3800 537.1500 1720.0000 ;
      RECT 527.4500 1719.3800 532.1500 1720.0000 ;
      RECT 522.4500 1719.3800 527.1500 1720.0000 ;
      RECT 517.4500 1719.3800 522.1500 1720.0000 ;
      RECT 512.4500 1719.3800 517.1500 1720.0000 ;
      RECT 507.4500 1719.3800 512.1500 1720.0000 ;
      RECT 502.4500 1719.3800 507.1500 1720.0000 ;
      RECT 497.4500 1719.3800 502.1500 1720.0000 ;
      RECT 492.4500 1719.3800 497.1500 1720.0000 ;
      RECT 487.4500 1719.3800 492.1500 1720.0000 ;
      RECT 482.4500 1719.3800 487.1500 1720.0000 ;
      RECT 477.4500 1719.3800 482.1500 1720.0000 ;
      RECT 472.4500 1719.3800 477.1500 1720.0000 ;
      RECT 467.4500 1719.3800 472.1500 1720.0000 ;
      RECT 462.4500 1719.3800 467.1500 1720.0000 ;
      RECT 457.4500 1719.3800 462.1500 1720.0000 ;
      RECT 452.4500 1719.3800 457.1500 1720.0000 ;
      RECT 447.4500 1719.3800 452.1500 1720.0000 ;
      RECT 442.4500 1719.3800 447.1500 1720.0000 ;
      RECT 437.4500 1719.3800 442.1500 1720.0000 ;
      RECT 432.4500 1719.3800 437.1500 1720.0000 ;
      RECT 427.4500 1719.3800 432.1500 1720.0000 ;
      RECT 422.4500 1719.3800 427.1500 1720.0000 ;
      RECT 417.4500 1719.3800 422.1500 1720.0000 ;
      RECT 412.4500 1719.3800 417.1500 1720.0000 ;
      RECT 407.4500 1719.3800 412.1500 1720.0000 ;
      RECT 402.4500 1719.3800 407.1500 1720.0000 ;
      RECT 397.4500 1719.3800 402.1500 1720.0000 ;
      RECT 392.4500 1719.3800 397.1500 1720.0000 ;
      RECT 387.4500 1719.3800 392.1500 1720.0000 ;
      RECT 382.4500 1719.3800 387.1500 1720.0000 ;
      RECT 377.4500 1719.3800 382.1500 1720.0000 ;
      RECT 372.4500 1719.3800 377.1500 1720.0000 ;
      RECT 367.4500 1719.3800 372.1500 1720.0000 ;
      RECT 362.4500 1719.3800 367.1500 1720.0000 ;
      RECT 357.4500 1719.3800 362.1500 1720.0000 ;
      RECT 352.4500 1719.3800 357.1500 1720.0000 ;
      RECT 347.4500 1719.3800 352.1500 1720.0000 ;
      RECT 342.4500 1719.3800 347.1500 1720.0000 ;
      RECT 337.4500 1719.3800 342.1500 1720.0000 ;
      RECT 332.4500 1719.3800 337.1500 1720.0000 ;
      RECT 327.4500 1719.3800 332.1500 1720.0000 ;
      RECT 322.4500 1719.3800 327.1500 1720.0000 ;
      RECT 317.4500 1719.3800 322.1500 1720.0000 ;
      RECT 312.4500 1719.3800 317.1500 1720.0000 ;
      RECT 307.4500 1719.3800 312.1500 1720.0000 ;
      RECT 302.4500 1719.3800 307.1500 1720.0000 ;
      RECT 297.4500 1719.3800 302.1500 1720.0000 ;
      RECT 292.4500 1719.3800 297.1500 1720.0000 ;
      RECT 287.4500 1719.3800 292.1500 1720.0000 ;
      RECT 282.4500 1719.3800 287.1500 1720.0000 ;
      RECT 277.4500 1719.3800 282.1500 1720.0000 ;
      RECT 272.4500 1719.3800 277.1500 1720.0000 ;
      RECT 267.4500 1719.3800 272.1500 1720.0000 ;
      RECT 262.4500 1719.3800 267.1500 1720.0000 ;
      RECT 257.4500 1719.3800 262.1500 1720.0000 ;
      RECT 252.4500 1719.3800 257.1500 1720.0000 ;
      RECT 247.4500 1719.3800 252.1500 1720.0000 ;
      RECT 242.4500 1719.3800 247.1500 1720.0000 ;
      RECT 237.4500 1719.3800 242.1500 1720.0000 ;
      RECT 232.4500 1719.3800 237.1500 1720.0000 ;
      RECT 0.0000 1719.3800 232.1500 1720.0000 ;
      RECT 0.0000 0.6200 1260.0000 1719.3800 ;
      RECT 1000.2500 0.0000 1260.0000 0.6200 ;
      RECT 995.2500 0.0000 999.9500 0.6200 ;
      RECT 990.2500 0.0000 994.9500 0.6200 ;
      RECT 985.2500 0.0000 989.9500 0.6200 ;
      RECT 980.2500 0.0000 984.9500 0.6200 ;
      RECT 975.2500 0.0000 979.9500 0.6200 ;
      RECT 970.2500 0.0000 974.9500 0.6200 ;
      RECT 965.2500 0.0000 969.9500 0.6200 ;
      RECT 960.2500 0.0000 964.9500 0.6200 ;
      RECT 955.2500 0.0000 959.9500 0.6200 ;
      RECT 950.2500 0.0000 954.9500 0.6200 ;
      RECT 945.2500 0.0000 949.9500 0.6200 ;
      RECT 940.2500 0.0000 944.9500 0.6200 ;
      RECT 935.2500 0.0000 939.9500 0.6200 ;
      RECT 930.2500 0.0000 934.9500 0.6200 ;
      RECT 925.2500 0.0000 929.9500 0.6200 ;
      RECT 920.2500 0.0000 924.9500 0.6200 ;
      RECT 915.2500 0.0000 919.9500 0.6200 ;
      RECT 910.2500 0.0000 914.9500 0.6200 ;
      RECT 905.2500 0.0000 909.9500 0.6200 ;
      RECT 900.2500 0.0000 904.9500 0.6200 ;
      RECT 895.2500 0.0000 899.9500 0.6200 ;
      RECT 890.2500 0.0000 894.9500 0.6200 ;
      RECT 885.2500 0.0000 889.9500 0.6200 ;
      RECT 880.2500 0.0000 884.9500 0.6200 ;
      RECT 875.2500 0.0000 879.9500 0.6200 ;
      RECT 870.2500 0.0000 874.9500 0.6200 ;
      RECT 865.2500 0.0000 869.9500 0.6200 ;
      RECT 860.2500 0.0000 864.9500 0.6200 ;
      RECT 855.2500 0.0000 859.9500 0.6200 ;
      RECT 850.2500 0.0000 854.9500 0.6200 ;
      RECT 845.2500 0.0000 849.9500 0.6200 ;
      RECT 840.2500 0.0000 844.9500 0.6200 ;
      RECT 835.2500 0.0000 839.9500 0.6200 ;
      RECT 830.2500 0.0000 834.9500 0.6200 ;
      RECT 825.2500 0.0000 829.9500 0.6200 ;
      RECT 820.2500 0.0000 824.9500 0.6200 ;
      RECT 815.2500 0.0000 819.9500 0.6200 ;
      RECT 810.2500 0.0000 814.9500 0.6200 ;
      RECT 805.2500 0.0000 809.9500 0.6200 ;
      RECT 800.2500 0.0000 804.9500 0.6200 ;
      RECT 795.2500 0.0000 799.9500 0.6200 ;
      RECT 790.2500 0.0000 794.9500 0.6200 ;
      RECT 785.2500 0.0000 789.9500 0.6200 ;
      RECT 780.2500 0.0000 784.9500 0.6200 ;
      RECT 775.2500 0.0000 779.9500 0.6200 ;
      RECT 770.2500 0.0000 774.9500 0.6200 ;
      RECT 765.2500 0.0000 769.9500 0.6200 ;
      RECT 760.2500 0.0000 764.9500 0.6200 ;
      RECT 755.2500 0.0000 759.9500 0.6200 ;
      RECT 750.2500 0.0000 754.9500 0.6200 ;
      RECT 745.2500 0.0000 749.9500 0.6200 ;
      RECT 740.2500 0.0000 744.9500 0.6200 ;
      RECT 735.2500 0.0000 739.9500 0.6200 ;
      RECT 730.2500 0.0000 734.9500 0.6200 ;
      RECT 725.2500 0.0000 729.9500 0.6200 ;
      RECT 720.2500 0.0000 724.9500 0.6200 ;
      RECT 715.2500 0.0000 719.9500 0.6200 ;
      RECT 710.2500 0.0000 714.9500 0.6200 ;
      RECT 705.2500 0.0000 709.9500 0.6200 ;
      RECT 700.2500 0.0000 704.9500 0.6200 ;
      RECT 695.2500 0.0000 699.9500 0.6200 ;
      RECT 690.2500 0.0000 694.9500 0.6200 ;
      RECT 685.2500 0.0000 689.9500 0.6200 ;
      RECT 680.2500 0.0000 684.9500 0.6200 ;
      RECT 675.2500 0.0000 679.9500 0.6200 ;
      RECT 670.2500 0.0000 674.9500 0.6200 ;
      RECT 665.2500 0.0000 669.9500 0.6200 ;
      RECT 660.2500 0.0000 664.9500 0.6200 ;
      RECT 655.2500 0.0000 659.9500 0.6200 ;
      RECT 650.2500 0.0000 654.9500 0.6200 ;
      RECT 645.2500 0.0000 649.9500 0.6200 ;
      RECT 640.2500 0.0000 644.9500 0.6200 ;
      RECT 635.2500 0.0000 639.9500 0.6200 ;
      RECT 630.2500 0.0000 634.9500 0.6200 ;
      RECT 625.2500 0.0000 629.9500 0.6200 ;
      RECT 620.2500 0.0000 624.9500 0.6200 ;
      RECT 615.2500 0.0000 619.9500 0.6200 ;
      RECT 610.2500 0.0000 614.9500 0.6200 ;
      RECT 605.2500 0.0000 609.9500 0.6200 ;
      RECT 600.2500 0.0000 604.9500 0.6200 ;
      RECT 595.2500 0.0000 599.9500 0.6200 ;
      RECT 590.2500 0.0000 594.9500 0.6200 ;
      RECT 585.2500 0.0000 589.9500 0.6200 ;
      RECT 580.2500 0.0000 584.9500 0.6200 ;
      RECT 575.2500 0.0000 579.9500 0.6200 ;
      RECT 570.2500 0.0000 574.9500 0.6200 ;
      RECT 565.2500 0.0000 569.9500 0.6200 ;
      RECT 560.2500 0.0000 564.9500 0.6200 ;
      RECT 555.2500 0.0000 559.9500 0.6200 ;
      RECT 550.2500 0.0000 554.9500 0.6200 ;
      RECT 545.2500 0.0000 549.9500 0.6200 ;
      RECT 540.2500 0.0000 544.9500 0.6200 ;
      RECT 535.2500 0.0000 539.9500 0.6200 ;
      RECT 530.2500 0.0000 534.9500 0.6200 ;
      RECT 525.2500 0.0000 529.9500 0.6200 ;
      RECT 520.2500 0.0000 524.9500 0.6200 ;
      RECT 515.2500 0.0000 519.9500 0.6200 ;
      RECT 510.2500 0.0000 514.9500 0.6200 ;
      RECT 505.2500 0.0000 509.9500 0.6200 ;
      RECT 500.2500 0.0000 504.9500 0.6200 ;
      RECT 495.2500 0.0000 499.9500 0.6200 ;
      RECT 490.2500 0.0000 494.9500 0.6200 ;
      RECT 485.2500 0.0000 489.9500 0.6200 ;
      RECT 480.2500 0.0000 484.9500 0.6200 ;
      RECT 475.2500 0.0000 479.9500 0.6200 ;
      RECT 470.2500 0.0000 474.9500 0.6200 ;
      RECT 465.2500 0.0000 469.9500 0.6200 ;
      RECT 460.2500 0.0000 464.9500 0.6200 ;
      RECT 455.2500 0.0000 459.9500 0.6200 ;
      RECT 450.2500 0.0000 454.9500 0.6200 ;
      RECT 445.2500 0.0000 449.9500 0.6200 ;
      RECT 440.2500 0.0000 444.9500 0.6200 ;
      RECT 435.2500 0.0000 439.9500 0.6200 ;
      RECT 430.2500 0.0000 434.9500 0.6200 ;
      RECT 425.2500 0.0000 429.9500 0.6200 ;
      RECT 420.2500 0.0000 424.9500 0.6200 ;
      RECT 415.2500 0.0000 419.9500 0.6200 ;
      RECT 410.2500 0.0000 414.9500 0.6200 ;
      RECT 405.2500 0.0000 409.9500 0.6200 ;
      RECT 400.2500 0.0000 404.9500 0.6200 ;
      RECT 395.2500 0.0000 399.9500 0.6200 ;
      RECT 390.2500 0.0000 394.9500 0.6200 ;
      RECT 385.2500 0.0000 389.9500 0.6200 ;
      RECT 380.2500 0.0000 384.9500 0.6200 ;
      RECT 375.2500 0.0000 379.9500 0.6200 ;
      RECT 370.2500 0.0000 374.9500 0.6200 ;
      RECT 365.2500 0.0000 369.9500 0.6200 ;
      RECT 360.2500 0.0000 364.9500 0.6200 ;
      RECT 355.2500 0.0000 359.9500 0.6200 ;
      RECT 350.2500 0.0000 354.9500 0.6200 ;
      RECT 345.2500 0.0000 349.9500 0.6200 ;
      RECT 340.2500 0.0000 344.9500 0.6200 ;
      RECT 335.2500 0.0000 339.9500 0.6200 ;
      RECT 330.2500 0.0000 334.9500 0.6200 ;
      RECT 325.2500 0.0000 329.9500 0.6200 ;
      RECT 320.2500 0.0000 324.9500 0.6200 ;
      RECT 315.2500 0.0000 319.9500 0.6200 ;
      RECT 310.2500 0.0000 314.9500 0.6200 ;
      RECT 305.2500 0.0000 309.9500 0.6200 ;
      RECT 300.2500 0.0000 304.9500 0.6200 ;
      RECT 295.2500 0.0000 299.9500 0.6200 ;
      RECT 290.2500 0.0000 294.9500 0.6200 ;
      RECT 285.2500 0.0000 289.9500 0.6200 ;
      RECT 280.2500 0.0000 284.9500 0.6200 ;
      RECT 275.2500 0.0000 279.9500 0.6200 ;
      RECT 270.2500 0.0000 274.9500 0.6200 ;
      RECT 265.2500 0.0000 269.9500 0.6200 ;
      RECT 260.2500 0.0000 264.9500 0.6200 ;
      RECT 0.0000 0.0000 259.9500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 980.3500 1260.0000 1720.0000 ;
      RECT 0.6200 980.0500 1260.0000 980.3500 ;
      RECT 0.0000 975.3500 1260.0000 980.0500 ;
      RECT 0.6200 975.0500 1260.0000 975.3500 ;
      RECT 0.0000 970.3500 1260.0000 975.0500 ;
      RECT 0.6200 970.0500 1260.0000 970.3500 ;
      RECT 0.0000 965.3500 1260.0000 970.0500 ;
      RECT 0.6200 965.0500 1260.0000 965.3500 ;
      RECT 0.0000 960.3500 1260.0000 965.0500 ;
      RECT 0.6200 960.0500 1260.0000 960.3500 ;
      RECT 0.0000 955.3500 1260.0000 960.0500 ;
      RECT 0.6200 955.0500 1260.0000 955.3500 ;
      RECT 0.0000 950.3500 1260.0000 955.0500 ;
      RECT 0.6200 950.0500 1260.0000 950.3500 ;
      RECT 0.0000 945.3500 1260.0000 950.0500 ;
      RECT 0.6200 945.0500 1260.0000 945.3500 ;
      RECT 0.0000 940.3500 1260.0000 945.0500 ;
      RECT 0.6200 940.0500 1260.0000 940.3500 ;
      RECT 0.0000 935.3500 1260.0000 940.0500 ;
      RECT 0.6200 935.0500 1260.0000 935.3500 ;
      RECT 0.0000 930.3500 1260.0000 935.0500 ;
      RECT 0.6200 930.0500 1260.0000 930.3500 ;
      RECT 0.0000 925.3500 1260.0000 930.0500 ;
      RECT 0.6200 925.0500 1260.0000 925.3500 ;
      RECT 0.0000 920.3500 1260.0000 925.0500 ;
      RECT 0.6200 920.0500 1260.0000 920.3500 ;
      RECT 0.0000 915.3500 1260.0000 920.0500 ;
      RECT 0.6200 915.0500 1260.0000 915.3500 ;
      RECT 0.0000 910.3500 1260.0000 915.0500 ;
      RECT 0.6200 910.0500 1260.0000 910.3500 ;
      RECT 0.0000 905.3500 1260.0000 910.0500 ;
      RECT 0.6200 905.0500 1260.0000 905.3500 ;
      RECT 0.0000 900.3500 1260.0000 905.0500 ;
      RECT 0.6200 900.0500 1260.0000 900.3500 ;
      RECT 0.0000 895.3500 1260.0000 900.0500 ;
      RECT 0.6200 895.0500 1260.0000 895.3500 ;
      RECT 0.0000 890.3500 1260.0000 895.0500 ;
      RECT 0.6200 890.0500 1260.0000 890.3500 ;
      RECT 0.0000 885.3500 1260.0000 890.0500 ;
      RECT 0.6200 885.0500 1260.0000 885.3500 ;
      RECT 0.0000 880.3500 1260.0000 885.0500 ;
      RECT 0.6200 880.0500 1260.0000 880.3500 ;
      RECT 0.0000 875.3500 1260.0000 880.0500 ;
      RECT 0.6200 875.0500 1260.0000 875.3500 ;
      RECT 0.0000 870.3500 1260.0000 875.0500 ;
      RECT 0.6200 870.0500 1260.0000 870.3500 ;
      RECT 0.0000 865.3500 1260.0000 870.0500 ;
      RECT 0.6200 865.0500 1260.0000 865.3500 ;
      RECT 0.0000 860.3500 1260.0000 865.0500 ;
      RECT 0.6200 860.0500 1260.0000 860.3500 ;
      RECT 0.0000 855.3500 1260.0000 860.0500 ;
      RECT 0.6200 855.0500 1260.0000 855.3500 ;
      RECT 0.0000 850.3500 1260.0000 855.0500 ;
      RECT 0.6200 850.0500 1260.0000 850.3500 ;
      RECT 0.0000 845.3500 1260.0000 850.0500 ;
      RECT 0.6200 845.0500 1260.0000 845.3500 ;
      RECT 0.0000 840.3500 1260.0000 845.0500 ;
      RECT 0.6200 840.0500 1260.0000 840.3500 ;
      RECT 0.0000 835.3500 1260.0000 840.0500 ;
      RECT 0.6200 835.0500 1260.0000 835.3500 ;
      RECT 0.0000 830.3500 1260.0000 835.0500 ;
      RECT 0.6200 830.0500 1260.0000 830.3500 ;
      RECT 0.0000 825.3500 1260.0000 830.0500 ;
      RECT 0.6200 825.0500 1260.0000 825.3500 ;
      RECT 0.0000 820.3500 1260.0000 825.0500 ;
      RECT 0.6200 820.0500 1260.0000 820.3500 ;
      RECT 0.0000 815.3500 1260.0000 820.0500 ;
      RECT 0.6200 815.0500 1260.0000 815.3500 ;
      RECT 0.0000 810.3500 1260.0000 815.0500 ;
      RECT 0.6200 810.0500 1260.0000 810.3500 ;
      RECT 0.0000 805.3500 1260.0000 810.0500 ;
      RECT 0.6200 805.0500 1260.0000 805.3500 ;
      RECT 0.0000 800.3500 1260.0000 805.0500 ;
      RECT 0.6200 800.0500 1260.0000 800.3500 ;
      RECT 0.0000 795.3500 1260.0000 800.0500 ;
      RECT 0.6200 795.0500 1260.0000 795.3500 ;
      RECT 0.0000 790.3500 1260.0000 795.0500 ;
      RECT 0.6200 790.0500 1260.0000 790.3500 ;
      RECT 0.0000 785.3500 1260.0000 790.0500 ;
      RECT 0.6200 785.0500 1260.0000 785.3500 ;
      RECT 0.0000 780.3500 1260.0000 785.0500 ;
      RECT 0.6200 780.0500 1260.0000 780.3500 ;
      RECT 0.0000 775.3500 1260.0000 780.0500 ;
      RECT 0.6200 775.0500 1260.0000 775.3500 ;
      RECT 0.0000 770.3500 1260.0000 775.0500 ;
      RECT 0.6200 770.0500 1260.0000 770.3500 ;
      RECT 0.0000 765.3500 1260.0000 770.0500 ;
      RECT 0.6200 765.0500 1260.0000 765.3500 ;
      RECT 0.0000 760.3500 1260.0000 765.0500 ;
      RECT 0.6200 760.0500 1260.0000 760.3500 ;
      RECT 0.0000 755.3500 1260.0000 760.0500 ;
      RECT 0.6200 755.0500 1260.0000 755.3500 ;
      RECT 0.0000 750.3500 1260.0000 755.0500 ;
      RECT 0.6200 750.0500 1260.0000 750.3500 ;
      RECT 0.0000 745.3500 1260.0000 750.0500 ;
      RECT 0.6200 745.0500 1260.0000 745.3500 ;
      RECT 0.0000 740.3500 1260.0000 745.0500 ;
      RECT 0.6200 740.0500 1260.0000 740.3500 ;
      RECT 0.0000 0.0000 1260.0000 740.0500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1260.0000 1720.0000 ;
  END
END core

END LIBRARY
