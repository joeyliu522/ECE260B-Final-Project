##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Mon Mar  3 16:56:45 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 695.6000 BY 695.0000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.3500 0.6000 55.4500 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 530.6500 0.0000 530.7500 0.5200 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 528.6500 0.0000 528.7500 0.5200 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 526.6500 0.0000 526.7500 0.5200 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 524.6500 0.0000 524.7500 0.5200 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 522.6500 0.0000 522.7500 0.5200 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 520.6500 0.0000 520.7500 0.5200 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 518.6500 0.0000 518.7500 0.5200 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 516.6500 0.0000 516.7500 0.5200 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 514.6500 0.0000 514.7500 0.5200 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 512.6500 0.0000 512.7500 0.5200 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.6500 0.0000 510.7500 0.5200 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 508.6500 0.0000 508.7500 0.5200 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 506.6500 0.0000 506.7500 0.5200 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 504.6500 0.0000 504.7500 0.5200 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 502.6500 0.0000 502.7500 0.5200 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.6500 0.0000 500.7500 0.5200 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 498.6500 0.0000 498.7500 0.5200 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 496.6500 0.0000 496.7500 0.5200 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 494.6500 0.0000 494.7500 0.5200 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.6500 0.0000 492.7500 0.5200 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 490.6500 0.0000 490.7500 0.5200 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 488.6500 0.0000 488.7500 0.5200 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 486.6500 0.0000 486.7500 0.5200 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 484.6500 0.0000 484.7500 0.5200 ;
    END
  END sum_out[0]
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 635.3500 0.6000 635.4500 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 631.3500 0.6000 631.4500 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 627.3500 0.6000 627.4500 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 623.3500 0.6000 623.4500 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 619.3500 0.6000 619.4500 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 615.3500 0.6000 615.4500 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 611.3500 0.6000 611.4500 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 607.3500 0.6000 607.4500 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 603.3500 0.6000 603.4500 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 599.3500 0.6000 599.4500 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 595.3500 0.6000 595.4500 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 591.3500 0.6000 591.4500 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 587.3500 0.6000 587.4500 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 583.3500 0.6000 583.4500 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 579.3500 0.6000 579.4500 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 575.3500 0.6000 575.4500 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 571.3500 0.6000 571.4500 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 567.3500 0.6000 567.4500 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 563.3500 0.6000 563.4500 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 559.3500 0.6000 559.4500 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 555.3500 0.6000 555.4500 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 551.3500 0.6000 551.4500 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 547.3500 0.6000 547.4500 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 543.3500 0.6000 543.4500 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 539.3500 0.6000 539.4500 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 535.3500 0.6000 535.4500 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 531.3500 0.6000 531.4500 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 527.3500 0.6000 527.4500 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 523.3500 0.6000 523.4500 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 519.3500 0.6000 519.4500 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 515.3500 0.6000 515.4500 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 511.3500 0.6000 511.4500 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 507.3500 0.6000 507.4500 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 503.3500 0.6000 503.4500 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 499.3500 0.6000 499.4500 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 495.3500 0.6000 495.4500 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 491.3500 0.6000 491.4500 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 487.3500 0.6000 487.4500 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 483.3500 0.6000 483.4500 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 479.3500 0.6000 479.4500 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 475.3500 0.6000 475.4500 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 471.3500 0.6000 471.4500 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 467.3500 0.6000 467.4500 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 463.3500 0.6000 463.4500 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 459.3500 0.6000 459.4500 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 455.3500 0.6000 455.4500 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 451.3500 0.6000 451.4500 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 447.3500 0.6000 447.4500 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 443.3500 0.6000 443.4500 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 439.3500 0.6000 439.4500 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 435.3500 0.6000 435.4500 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 431.3500 0.6000 431.4500 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 427.3500 0.6000 427.4500 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 423.3500 0.6000 423.4500 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 419.3500 0.6000 419.4500 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 415.3500 0.6000 415.4500 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 411.3500 0.6000 411.4500 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 407.3500 0.6000 407.4500 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 403.3500 0.6000 403.4500 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 399.3500 0.6000 399.4500 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 395.3500 0.6000 395.4500 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 391.3500 0.6000 391.4500 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 387.3500 0.6000 387.4500 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 383.3500 0.6000 383.4500 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 379.3500 0.6000 379.4500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 375.3500 0.6000 375.4500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 371.3500 0.6000 371.4500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 367.3500 0.6000 367.4500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 363.3500 0.6000 363.4500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 359.3500 0.6000 359.4500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 355.3500 0.6000 355.4500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 351.3500 0.6000 351.4500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 347.3500 0.6000 347.4500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 343.3500 0.6000 343.4500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 339.3500 0.6000 339.4500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 335.3500 0.6000 335.4500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 331.3500 0.6000 331.4500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 327.3500 0.6000 327.4500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 323.3500 0.6000 323.4500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 319.3500 0.6000 319.4500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 315.3500 0.6000 315.4500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 311.3500 0.6000 311.4500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 307.3500 0.6000 307.4500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 303.3500 0.6000 303.4500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 299.3500 0.6000 299.4500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 295.3500 0.6000 295.4500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 291.3500 0.6000 291.4500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 287.3500 0.6000 287.4500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 283.3500 0.6000 283.4500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 279.3500 0.6000 279.4500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 275.3500 0.6000 275.4500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 271.3500 0.6000 271.4500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 267.3500 0.6000 267.4500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 263.3500 0.6000 263.4500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 259.3500 0.6000 259.4500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 255.3500 0.6000 255.4500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 251.3500 0.6000 251.4500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 247.3500 0.6000 247.4500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 243.3500 0.6000 243.4500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 239.3500 0.6000 239.4500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 235.3500 0.6000 235.4500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 231.3500 0.6000 231.4500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 227.3500 0.6000 227.4500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 223.3500 0.6000 223.4500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 219.3500 0.6000 219.4500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.3500 0.6000 215.4500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.3500 0.6000 211.4500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 207.3500 0.6000 207.4500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 203.3500 0.6000 203.4500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 199.3500 0.6000 199.4500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.3500 0.6000 195.4500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 191.3500 0.6000 191.4500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 187.3500 0.6000 187.4500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 183.3500 0.6000 183.4500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 179.3500 0.6000 179.4500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 175.3500 0.6000 175.4500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 171.3500 0.6000 171.4500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 167.3500 0.6000 167.4500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 163.3500 0.6000 163.4500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 159.3500 0.6000 159.4500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 155.3500 0.6000 155.4500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 151.3500 0.6000 151.4500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 147.3500 0.6000 147.4500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 143.3500 0.6000 143.4500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 139.3500 0.6000 139.4500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 135.3500 0.6000 135.4500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 131.3500 0.6000 131.4500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 127.3500 0.6000 127.4500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 482.6500 0.0000 482.7500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 480.6500 0.0000 480.7500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.6500 0.0000 478.7500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 476.6500 0.0000 476.7500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 474.6500 0.0000 474.7500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 472.6500 0.0000 472.7500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.6500 0.0000 470.7500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 468.6500 0.0000 468.7500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 466.6500 0.0000 466.7500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.6500 0.0000 464.7500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 462.6500 0.0000 462.7500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.6500 0.0000 460.7500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.6500 0.0000 458.7500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.6500 0.0000 456.7500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.6500 0.0000 454.7500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.6500 0.0000 452.7500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.6500 0.0000 450.7500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.6500 0.0000 448.7500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.6500 0.0000 446.7500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.6500 0.0000 444.7500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.6500 0.0000 442.7500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.6500 0.0000 440.7500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.6500 0.0000 438.7500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.6500 0.0000 436.7500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.6500 0.0000 434.7500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.6500 0.0000 432.7500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.6500 0.0000 430.7500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.6500 0.0000 428.7500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.6500 0.0000 426.7500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.6500 0.0000 424.7500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.6500 0.0000 422.7500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.6500 0.0000 420.7500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.6500 0.0000 418.7500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.6500 0.0000 416.7500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.6500 0.0000 414.7500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.6500 0.0000 412.7500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.6500 0.0000 410.7500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.6500 0.0000 408.7500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.6500 0.0000 406.7500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.6500 0.0000 404.7500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.6500 0.0000 402.7500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.6500 0.0000 400.7500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.6500 0.0000 398.7500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.6500 0.0000 396.7500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.6500 0.0000 394.7500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.6500 0.0000 392.7500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.6500 0.0000 390.7500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.6500 0.0000 388.7500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.6500 0.0000 386.7500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.6500 0.0000 384.7500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.6500 0.0000 382.7500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.6500 0.0000 380.7500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.6500 0.0000 378.7500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.6500 0.0000 376.7500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.6500 0.0000 374.7500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.6500 0.0000 372.7500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.6500 0.0000 370.7500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.6500 0.0000 368.7500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.6500 0.0000 366.7500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.6500 0.0000 364.7500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.6500 0.0000 362.7500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.6500 0.0000 360.7500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.6500 0.0000 358.7500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.6500 0.0000 356.7500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.6500 0.0000 354.7500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.6500 0.0000 352.7500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.6500 0.0000 350.7500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.6500 0.0000 348.7500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.6500 0.0000 346.7500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.6500 0.0000 344.7500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.6500 0.0000 342.7500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.6500 0.0000 340.7500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.6500 0.0000 338.7500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.6500 0.0000 336.7500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.6500 0.0000 334.7500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.6500 0.0000 332.7500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.6500 0.0000 330.7500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.6500 0.0000 328.7500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.6500 0.0000 326.7500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.6500 0.0000 324.7500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.6500 0.0000 322.7500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.6500 0.0000 320.7500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.6500 0.0000 318.7500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.6500 0.0000 316.7500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.6500 0.0000 314.7500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.6500 0.0000 312.7500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.6500 0.0000 310.7500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.6500 0.0000 308.7500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.6500 0.0000 306.7500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.6500 0.0000 304.7500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.6500 0.0000 302.7500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.6500 0.0000 300.7500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.6500 0.0000 298.7500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.6500 0.0000 296.7500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.6500 0.0000 294.7500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.6500 0.0000 292.7500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.6500 0.0000 290.7500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.6500 0.0000 288.7500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.6500 0.0000 286.7500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.6500 0.0000 284.7500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.6500 0.0000 282.7500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.6500 0.0000 280.7500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.6500 0.0000 278.7500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.6500 0.0000 276.7500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.6500 0.0000 274.7500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.6500 0.0000 272.7500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.6500 0.0000 270.7500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.6500 0.0000 268.7500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.6500 0.0000 266.7500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.6500 0.0000 264.7500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.6500 0.0000 262.7500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.6500 0.0000 260.7500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.6500 0.0000 258.7500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.6500 0.0000 256.7500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.6500 0.0000 254.7500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.6500 0.0000 252.7500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.6500 0.0000 250.7500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.6500 0.0000 248.7500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.6500 0.0000 246.7500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.6500 0.0000 244.7500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.6500 0.0000 242.7500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.6500 0.0000 240.7500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.6500 0.0000 238.7500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.6500 0.0000 236.7500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.6500 0.0000 234.7500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.6500 0.0000 232.7500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.6500 0.0000 230.7500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.6500 0.0000 228.7500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.6500 0.0000 226.7500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.6500 0.0000 224.7500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.6500 0.0000 222.7500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.6500 0.0000 220.7500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.6500 0.0000 218.7500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.6500 0.0000 216.7500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.6500 0.0000 214.7500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.6500 0.0000 212.7500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.6500 0.0000 210.7500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.6500 0.0000 208.7500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.6500 0.0000 206.7500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.6500 0.0000 204.7500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.6500 0.0000 202.7500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.6500 0.0000 200.7500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.6500 0.0000 198.7500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.6500 0.0000 196.7500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.6500 0.0000 194.7500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.6500 0.0000 192.7500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.6500 0.0000 190.7500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.6500 0.0000 188.7500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.6500 0.0000 186.7500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.6500 0.0000 184.7500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.6500 0.0000 182.7500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.6500 0.0000 180.7500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.6500 0.0000 178.7500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.6500 0.0000 176.7500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.6500 0.0000 174.7500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.6500 0.0000 172.7500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.6500 0.0000 170.7500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.6500 0.0000 168.7500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.6500 0.0000 166.7500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.6500 0.0000 164.7500 0.5200 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 123.3500 0.6000 123.4500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 119.3500 0.6000 119.4500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 115.3500 0.6000 115.4500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 111.3500 0.6000 111.4500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 107.3500 0.6000 107.4500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 103.3500 0.6000 103.4500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 99.3500 0.6000 99.4500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 95.3500 0.6000 95.4500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 91.3500 0.6000 91.4500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 87.3500 0.6000 87.4500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 83.3500 0.6000 83.4500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 79.3500 0.6000 79.4500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 75.3500 0.6000 75.4500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 71.3500 0.6000 71.4500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 67.3500 0.6000 67.4500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.3500 0.6000 63.4500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.3500 0.6000 59.4500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 639.3500 0.6000 639.4500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.6200 695.6000 695.0000 ;
      RECT 530.8500 0.0000 695.6000 0.6200 ;
      RECT 528.8500 0.0000 530.5500 0.6200 ;
      RECT 526.8500 0.0000 528.5500 0.6200 ;
      RECT 524.8500 0.0000 526.5500 0.6200 ;
      RECT 522.8500 0.0000 524.5500 0.6200 ;
      RECT 520.8500 0.0000 522.5500 0.6200 ;
      RECT 518.8500 0.0000 520.5500 0.6200 ;
      RECT 516.8500 0.0000 518.5500 0.6200 ;
      RECT 514.8500 0.0000 516.5500 0.6200 ;
      RECT 512.8500 0.0000 514.5500 0.6200 ;
      RECT 510.8500 0.0000 512.5500 0.6200 ;
      RECT 508.8500 0.0000 510.5500 0.6200 ;
      RECT 506.8500 0.0000 508.5500 0.6200 ;
      RECT 504.8500 0.0000 506.5500 0.6200 ;
      RECT 502.8500 0.0000 504.5500 0.6200 ;
      RECT 500.8500 0.0000 502.5500 0.6200 ;
      RECT 498.8500 0.0000 500.5500 0.6200 ;
      RECT 496.8500 0.0000 498.5500 0.6200 ;
      RECT 494.8500 0.0000 496.5500 0.6200 ;
      RECT 492.8500 0.0000 494.5500 0.6200 ;
      RECT 490.8500 0.0000 492.5500 0.6200 ;
      RECT 488.8500 0.0000 490.5500 0.6200 ;
      RECT 486.8500 0.0000 488.5500 0.6200 ;
      RECT 484.8500 0.0000 486.5500 0.6200 ;
      RECT 482.8500 0.0000 484.5500 0.6200 ;
      RECT 480.8500 0.0000 482.5500 0.6200 ;
      RECT 478.8500 0.0000 480.5500 0.6200 ;
      RECT 476.8500 0.0000 478.5500 0.6200 ;
      RECT 474.8500 0.0000 476.5500 0.6200 ;
      RECT 472.8500 0.0000 474.5500 0.6200 ;
      RECT 470.8500 0.0000 472.5500 0.6200 ;
      RECT 468.8500 0.0000 470.5500 0.6200 ;
      RECT 466.8500 0.0000 468.5500 0.6200 ;
      RECT 464.8500 0.0000 466.5500 0.6200 ;
      RECT 462.8500 0.0000 464.5500 0.6200 ;
      RECT 460.8500 0.0000 462.5500 0.6200 ;
      RECT 458.8500 0.0000 460.5500 0.6200 ;
      RECT 456.8500 0.0000 458.5500 0.6200 ;
      RECT 454.8500 0.0000 456.5500 0.6200 ;
      RECT 452.8500 0.0000 454.5500 0.6200 ;
      RECT 450.8500 0.0000 452.5500 0.6200 ;
      RECT 448.8500 0.0000 450.5500 0.6200 ;
      RECT 446.8500 0.0000 448.5500 0.6200 ;
      RECT 444.8500 0.0000 446.5500 0.6200 ;
      RECT 442.8500 0.0000 444.5500 0.6200 ;
      RECT 440.8500 0.0000 442.5500 0.6200 ;
      RECT 438.8500 0.0000 440.5500 0.6200 ;
      RECT 436.8500 0.0000 438.5500 0.6200 ;
      RECT 434.8500 0.0000 436.5500 0.6200 ;
      RECT 432.8500 0.0000 434.5500 0.6200 ;
      RECT 430.8500 0.0000 432.5500 0.6200 ;
      RECT 428.8500 0.0000 430.5500 0.6200 ;
      RECT 426.8500 0.0000 428.5500 0.6200 ;
      RECT 424.8500 0.0000 426.5500 0.6200 ;
      RECT 422.8500 0.0000 424.5500 0.6200 ;
      RECT 420.8500 0.0000 422.5500 0.6200 ;
      RECT 418.8500 0.0000 420.5500 0.6200 ;
      RECT 416.8500 0.0000 418.5500 0.6200 ;
      RECT 414.8500 0.0000 416.5500 0.6200 ;
      RECT 412.8500 0.0000 414.5500 0.6200 ;
      RECT 410.8500 0.0000 412.5500 0.6200 ;
      RECT 408.8500 0.0000 410.5500 0.6200 ;
      RECT 406.8500 0.0000 408.5500 0.6200 ;
      RECT 404.8500 0.0000 406.5500 0.6200 ;
      RECT 402.8500 0.0000 404.5500 0.6200 ;
      RECT 400.8500 0.0000 402.5500 0.6200 ;
      RECT 398.8500 0.0000 400.5500 0.6200 ;
      RECT 396.8500 0.0000 398.5500 0.6200 ;
      RECT 394.8500 0.0000 396.5500 0.6200 ;
      RECT 392.8500 0.0000 394.5500 0.6200 ;
      RECT 390.8500 0.0000 392.5500 0.6200 ;
      RECT 388.8500 0.0000 390.5500 0.6200 ;
      RECT 386.8500 0.0000 388.5500 0.6200 ;
      RECT 384.8500 0.0000 386.5500 0.6200 ;
      RECT 382.8500 0.0000 384.5500 0.6200 ;
      RECT 380.8500 0.0000 382.5500 0.6200 ;
      RECT 378.8500 0.0000 380.5500 0.6200 ;
      RECT 376.8500 0.0000 378.5500 0.6200 ;
      RECT 374.8500 0.0000 376.5500 0.6200 ;
      RECT 372.8500 0.0000 374.5500 0.6200 ;
      RECT 370.8500 0.0000 372.5500 0.6200 ;
      RECT 368.8500 0.0000 370.5500 0.6200 ;
      RECT 366.8500 0.0000 368.5500 0.6200 ;
      RECT 364.8500 0.0000 366.5500 0.6200 ;
      RECT 362.8500 0.0000 364.5500 0.6200 ;
      RECT 360.8500 0.0000 362.5500 0.6200 ;
      RECT 358.8500 0.0000 360.5500 0.6200 ;
      RECT 356.8500 0.0000 358.5500 0.6200 ;
      RECT 354.8500 0.0000 356.5500 0.6200 ;
      RECT 352.8500 0.0000 354.5500 0.6200 ;
      RECT 350.8500 0.0000 352.5500 0.6200 ;
      RECT 348.8500 0.0000 350.5500 0.6200 ;
      RECT 346.8500 0.0000 348.5500 0.6200 ;
      RECT 344.8500 0.0000 346.5500 0.6200 ;
      RECT 342.8500 0.0000 344.5500 0.6200 ;
      RECT 340.8500 0.0000 342.5500 0.6200 ;
      RECT 338.8500 0.0000 340.5500 0.6200 ;
      RECT 336.8500 0.0000 338.5500 0.6200 ;
      RECT 334.8500 0.0000 336.5500 0.6200 ;
      RECT 332.8500 0.0000 334.5500 0.6200 ;
      RECT 330.8500 0.0000 332.5500 0.6200 ;
      RECT 328.8500 0.0000 330.5500 0.6200 ;
      RECT 326.8500 0.0000 328.5500 0.6200 ;
      RECT 324.8500 0.0000 326.5500 0.6200 ;
      RECT 322.8500 0.0000 324.5500 0.6200 ;
      RECT 320.8500 0.0000 322.5500 0.6200 ;
      RECT 318.8500 0.0000 320.5500 0.6200 ;
      RECT 316.8500 0.0000 318.5500 0.6200 ;
      RECT 314.8500 0.0000 316.5500 0.6200 ;
      RECT 312.8500 0.0000 314.5500 0.6200 ;
      RECT 310.8500 0.0000 312.5500 0.6200 ;
      RECT 308.8500 0.0000 310.5500 0.6200 ;
      RECT 306.8500 0.0000 308.5500 0.6200 ;
      RECT 304.8500 0.0000 306.5500 0.6200 ;
      RECT 302.8500 0.0000 304.5500 0.6200 ;
      RECT 300.8500 0.0000 302.5500 0.6200 ;
      RECT 298.8500 0.0000 300.5500 0.6200 ;
      RECT 296.8500 0.0000 298.5500 0.6200 ;
      RECT 294.8500 0.0000 296.5500 0.6200 ;
      RECT 292.8500 0.0000 294.5500 0.6200 ;
      RECT 290.8500 0.0000 292.5500 0.6200 ;
      RECT 288.8500 0.0000 290.5500 0.6200 ;
      RECT 286.8500 0.0000 288.5500 0.6200 ;
      RECT 284.8500 0.0000 286.5500 0.6200 ;
      RECT 282.8500 0.0000 284.5500 0.6200 ;
      RECT 280.8500 0.0000 282.5500 0.6200 ;
      RECT 278.8500 0.0000 280.5500 0.6200 ;
      RECT 276.8500 0.0000 278.5500 0.6200 ;
      RECT 274.8500 0.0000 276.5500 0.6200 ;
      RECT 272.8500 0.0000 274.5500 0.6200 ;
      RECT 270.8500 0.0000 272.5500 0.6200 ;
      RECT 268.8500 0.0000 270.5500 0.6200 ;
      RECT 266.8500 0.0000 268.5500 0.6200 ;
      RECT 264.8500 0.0000 266.5500 0.6200 ;
      RECT 262.8500 0.0000 264.5500 0.6200 ;
      RECT 260.8500 0.0000 262.5500 0.6200 ;
      RECT 258.8500 0.0000 260.5500 0.6200 ;
      RECT 256.8500 0.0000 258.5500 0.6200 ;
      RECT 254.8500 0.0000 256.5500 0.6200 ;
      RECT 252.8500 0.0000 254.5500 0.6200 ;
      RECT 250.8500 0.0000 252.5500 0.6200 ;
      RECT 248.8500 0.0000 250.5500 0.6200 ;
      RECT 246.8500 0.0000 248.5500 0.6200 ;
      RECT 244.8500 0.0000 246.5500 0.6200 ;
      RECT 242.8500 0.0000 244.5500 0.6200 ;
      RECT 240.8500 0.0000 242.5500 0.6200 ;
      RECT 238.8500 0.0000 240.5500 0.6200 ;
      RECT 236.8500 0.0000 238.5500 0.6200 ;
      RECT 234.8500 0.0000 236.5500 0.6200 ;
      RECT 232.8500 0.0000 234.5500 0.6200 ;
      RECT 230.8500 0.0000 232.5500 0.6200 ;
      RECT 228.8500 0.0000 230.5500 0.6200 ;
      RECT 226.8500 0.0000 228.5500 0.6200 ;
      RECT 224.8500 0.0000 226.5500 0.6200 ;
      RECT 222.8500 0.0000 224.5500 0.6200 ;
      RECT 220.8500 0.0000 222.5500 0.6200 ;
      RECT 218.8500 0.0000 220.5500 0.6200 ;
      RECT 216.8500 0.0000 218.5500 0.6200 ;
      RECT 214.8500 0.0000 216.5500 0.6200 ;
      RECT 212.8500 0.0000 214.5500 0.6200 ;
      RECT 210.8500 0.0000 212.5500 0.6200 ;
      RECT 208.8500 0.0000 210.5500 0.6200 ;
      RECT 206.8500 0.0000 208.5500 0.6200 ;
      RECT 204.8500 0.0000 206.5500 0.6200 ;
      RECT 202.8500 0.0000 204.5500 0.6200 ;
      RECT 200.8500 0.0000 202.5500 0.6200 ;
      RECT 198.8500 0.0000 200.5500 0.6200 ;
      RECT 196.8500 0.0000 198.5500 0.6200 ;
      RECT 194.8500 0.0000 196.5500 0.6200 ;
      RECT 192.8500 0.0000 194.5500 0.6200 ;
      RECT 190.8500 0.0000 192.5500 0.6200 ;
      RECT 188.8500 0.0000 190.5500 0.6200 ;
      RECT 186.8500 0.0000 188.5500 0.6200 ;
      RECT 184.8500 0.0000 186.5500 0.6200 ;
      RECT 182.8500 0.0000 184.5500 0.6200 ;
      RECT 180.8500 0.0000 182.5500 0.6200 ;
      RECT 178.8500 0.0000 180.5500 0.6200 ;
      RECT 176.8500 0.0000 178.5500 0.6200 ;
      RECT 174.8500 0.0000 176.5500 0.6200 ;
      RECT 172.8500 0.0000 174.5500 0.6200 ;
      RECT 170.8500 0.0000 172.5500 0.6200 ;
      RECT 168.8500 0.0000 170.5500 0.6200 ;
      RECT 166.8500 0.0000 168.5500 0.6200 ;
      RECT 164.8500 0.0000 166.5500 0.6200 ;
      RECT 0.0000 0.0000 164.5500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 639.5500 695.6000 695.0000 ;
      RECT 0.7000 639.2500 695.6000 639.5500 ;
      RECT 0.0000 635.5500 695.6000 639.2500 ;
      RECT 0.7000 635.2500 695.6000 635.5500 ;
      RECT 0.0000 631.5500 695.6000 635.2500 ;
      RECT 0.7000 631.2500 695.6000 631.5500 ;
      RECT 0.0000 627.5500 695.6000 631.2500 ;
      RECT 0.7000 627.2500 695.6000 627.5500 ;
      RECT 0.0000 623.5500 695.6000 627.2500 ;
      RECT 0.7000 623.2500 695.6000 623.5500 ;
      RECT 0.0000 619.5500 695.6000 623.2500 ;
      RECT 0.7000 619.2500 695.6000 619.5500 ;
      RECT 0.0000 615.5500 695.6000 619.2500 ;
      RECT 0.7000 615.2500 695.6000 615.5500 ;
      RECT 0.0000 611.5500 695.6000 615.2500 ;
      RECT 0.7000 611.2500 695.6000 611.5500 ;
      RECT 0.0000 607.5500 695.6000 611.2500 ;
      RECT 0.7000 607.2500 695.6000 607.5500 ;
      RECT 0.0000 603.5500 695.6000 607.2500 ;
      RECT 0.7000 603.2500 695.6000 603.5500 ;
      RECT 0.0000 599.5500 695.6000 603.2500 ;
      RECT 0.7000 599.2500 695.6000 599.5500 ;
      RECT 0.0000 595.5500 695.6000 599.2500 ;
      RECT 0.7000 595.2500 695.6000 595.5500 ;
      RECT 0.0000 591.5500 695.6000 595.2500 ;
      RECT 0.7000 591.2500 695.6000 591.5500 ;
      RECT 0.0000 587.5500 695.6000 591.2500 ;
      RECT 0.7000 587.2500 695.6000 587.5500 ;
      RECT 0.0000 583.5500 695.6000 587.2500 ;
      RECT 0.7000 583.2500 695.6000 583.5500 ;
      RECT 0.0000 579.5500 695.6000 583.2500 ;
      RECT 0.7000 579.2500 695.6000 579.5500 ;
      RECT 0.0000 575.5500 695.6000 579.2500 ;
      RECT 0.7000 575.2500 695.6000 575.5500 ;
      RECT 0.0000 571.5500 695.6000 575.2500 ;
      RECT 0.7000 571.2500 695.6000 571.5500 ;
      RECT 0.0000 567.5500 695.6000 571.2500 ;
      RECT 0.7000 567.2500 695.6000 567.5500 ;
      RECT 0.0000 563.5500 695.6000 567.2500 ;
      RECT 0.7000 563.2500 695.6000 563.5500 ;
      RECT 0.0000 559.5500 695.6000 563.2500 ;
      RECT 0.7000 559.2500 695.6000 559.5500 ;
      RECT 0.0000 555.5500 695.6000 559.2500 ;
      RECT 0.7000 555.2500 695.6000 555.5500 ;
      RECT 0.0000 551.5500 695.6000 555.2500 ;
      RECT 0.7000 551.2500 695.6000 551.5500 ;
      RECT 0.0000 547.5500 695.6000 551.2500 ;
      RECT 0.7000 547.2500 695.6000 547.5500 ;
      RECT 0.0000 543.5500 695.6000 547.2500 ;
      RECT 0.7000 543.2500 695.6000 543.5500 ;
      RECT 0.0000 539.5500 695.6000 543.2500 ;
      RECT 0.7000 539.2500 695.6000 539.5500 ;
      RECT 0.0000 535.5500 695.6000 539.2500 ;
      RECT 0.7000 535.2500 695.6000 535.5500 ;
      RECT 0.0000 531.5500 695.6000 535.2500 ;
      RECT 0.7000 531.2500 695.6000 531.5500 ;
      RECT 0.0000 527.5500 695.6000 531.2500 ;
      RECT 0.7000 527.2500 695.6000 527.5500 ;
      RECT 0.0000 523.5500 695.6000 527.2500 ;
      RECT 0.7000 523.2500 695.6000 523.5500 ;
      RECT 0.0000 519.5500 695.6000 523.2500 ;
      RECT 0.7000 519.2500 695.6000 519.5500 ;
      RECT 0.0000 515.5500 695.6000 519.2500 ;
      RECT 0.7000 515.2500 695.6000 515.5500 ;
      RECT 0.0000 511.5500 695.6000 515.2500 ;
      RECT 0.7000 511.2500 695.6000 511.5500 ;
      RECT 0.0000 507.5500 695.6000 511.2500 ;
      RECT 0.7000 507.2500 695.6000 507.5500 ;
      RECT 0.0000 503.5500 695.6000 507.2500 ;
      RECT 0.7000 503.2500 695.6000 503.5500 ;
      RECT 0.0000 499.5500 695.6000 503.2500 ;
      RECT 0.7000 499.2500 695.6000 499.5500 ;
      RECT 0.0000 495.5500 695.6000 499.2500 ;
      RECT 0.7000 495.2500 695.6000 495.5500 ;
      RECT 0.0000 491.5500 695.6000 495.2500 ;
      RECT 0.7000 491.2500 695.6000 491.5500 ;
      RECT 0.0000 487.5500 695.6000 491.2500 ;
      RECT 0.7000 487.2500 695.6000 487.5500 ;
      RECT 0.0000 483.5500 695.6000 487.2500 ;
      RECT 0.7000 483.2500 695.6000 483.5500 ;
      RECT 0.0000 479.5500 695.6000 483.2500 ;
      RECT 0.7000 479.2500 695.6000 479.5500 ;
      RECT 0.0000 475.5500 695.6000 479.2500 ;
      RECT 0.7000 475.2500 695.6000 475.5500 ;
      RECT 0.0000 471.5500 695.6000 475.2500 ;
      RECT 0.7000 471.2500 695.6000 471.5500 ;
      RECT 0.0000 467.5500 695.6000 471.2500 ;
      RECT 0.7000 467.2500 695.6000 467.5500 ;
      RECT 0.0000 463.5500 695.6000 467.2500 ;
      RECT 0.7000 463.2500 695.6000 463.5500 ;
      RECT 0.0000 459.5500 695.6000 463.2500 ;
      RECT 0.7000 459.2500 695.6000 459.5500 ;
      RECT 0.0000 455.5500 695.6000 459.2500 ;
      RECT 0.7000 455.2500 695.6000 455.5500 ;
      RECT 0.0000 451.5500 695.6000 455.2500 ;
      RECT 0.7000 451.2500 695.6000 451.5500 ;
      RECT 0.0000 447.5500 695.6000 451.2500 ;
      RECT 0.7000 447.2500 695.6000 447.5500 ;
      RECT 0.0000 443.5500 695.6000 447.2500 ;
      RECT 0.7000 443.2500 695.6000 443.5500 ;
      RECT 0.0000 439.5500 695.6000 443.2500 ;
      RECT 0.7000 439.2500 695.6000 439.5500 ;
      RECT 0.0000 435.5500 695.6000 439.2500 ;
      RECT 0.7000 435.2500 695.6000 435.5500 ;
      RECT 0.0000 431.5500 695.6000 435.2500 ;
      RECT 0.7000 431.2500 695.6000 431.5500 ;
      RECT 0.0000 427.5500 695.6000 431.2500 ;
      RECT 0.7000 427.2500 695.6000 427.5500 ;
      RECT 0.0000 423.5500 695.6000 427.2500 ;
      RECT 0.7000 423.2500 695.6000 423.5500 ;
      RECT 0.0000 419.5500 695.6000 423.2500 ;
      RECT 0.7000 419.2500 695.6000 419.5500 ;
      RECT 0.0000 415.5500 695.6000 419.2500 ;
      RECT 0.7000 415.2500 695.6000 415.5500 ;
      RECT 0.0000 411.5500 695.6000 415.2500 ;
      RECT 0.7000 411.2500 695.6000 411.5500 ;
      RECT 0.0000 407.5500 695.6000 411.2500 ;
      RECT 0.7000 407.2500 695.6000 407.5500 ;
      RECT 0.0000 403.5500 695.6000 407.2500 ;
      RECT 0.7000 403.2500 695.6000 403.5500 ;
      RECT 0.0000 399.5500 695.6000 403.2500 ;
      RECT 0.7000 399.2500 695.6000 399.5500 ;
      RECT 0.0000 395.5500 695.6000 399.2500 ;
      RECT 0.7000 395.2500 695.6000 395.5500 ;
      RECT 0.0000 391.5500 695.6000 395.2500 ;
      RECT 0.7000 391.2500 695.6000 391.5500 ;
      RECT 0.0000 387.5500 695.6000 391.2500 ;
      RECT 0.7000 387.2500 695.6000 387.5500 ;
      RECT 0.0000 383.5500 695.6000 387.2500 ;
      RECT 0.7000 383.2500 695.6000 383.5500 ;
      RECT 0.0000 379.5500 695.6000 383.2500 ;
      RECT 0.7000 379.2500 695.6000 379.5500 ;
      RECT 0.0000 375.5500 695.6000 379.2500 ;
      RECT 0.7000 375.2500 695.6000 375.5500 ;
      RECT 0.0000 371.5500 695.6000 375.2500 ;
      RECT 0.7000 371.2500 695.6000 371.5500 ;
      RECT 0.0000 367.5500 695.6000 371.2500 ;
      RECT 0.7000 367.2500 695.6000 367.5500 ;
      RECT 0.0000 363.5500 695.6000 367.2500 ;
      RECT 0.7000 363.2500 695.6000 363.5500 ;
      RECT 0.0000 359.5500 695.6000 363.2500 ;
      RECT 0.7000 359.2500 695.6000 359.5500 ;
      RECT 0.0000 355.5500 695.6000 359.2500 ;
      RECT 0.7000 355.2500 695.6000 355.5500 ;
      RECT 0.0000 351.5500 695.6000 355.2500 ;
      RECT 0.7000 351.2500 695.6000 351.5500 ;
      RECT 0.0000 347.5500 695.6000 351.2500 ;
      RECT 0.7000 347.2500 695.6000 347.5500 ;
      RECT 0.0000 343.5500 695.6000 347.2500 ;
      RECT 0.7000 343.2500 695.6000 343.5500 ;
      RECT 0.0000 339.5500 695.6000 343.2500 ;
      RECT 0.7000 339.2500 695.6000 339.5500 ;
      RECT 0.0000 335.5500 695.6000 339.2500 ;
      RECT 0.7000 335.2500 695.6000 335.5500 ;
      RECT 0.0000 331.5500 695.6000 335.2500 ;
      RECT 0.7000 331.2500 695.6000 331.5500 ;
      RECT 0.0000 327.5500 695.6000 331.2500 ;
      RECT 0.7000 327.2500 695.6000 327.5500 ;
      RECT 0.0000 323.5500 695.6000 327.2500 ;
      RECT 0.7000 323.2500 695.6000 323.5500 ;
      RECT 0.0000 319.5500 695.6000 323.2500 ;
      RECT 0.7000 319.2500 695.6000 319.5500 ;
      RECT 0.0000 315.5500 695.6000 319.2500 ;
      RECT 0.7000 315.2500 695.6000 315.5500 ;
      RECT 0.0000 311.5500 695.6000 315.2500 ;
      RECT 0.7000 311.2500 695.6000 311.5500 ;
      RECT 0.0000 307.5500 695.6000 311.2500 ;
      RECT 0.7000 307.2500 695.6000 307.5500 ;
      RECT 0.0000 303.5500 695.6000 307.2500 ;
      RECT 0.7000 303.2500 695.6000 303.5500 ;
      RECT 0.0000 299.5500 695.6000 303.2500 ;
      RECT 0.7000 299.2500 695.6000 299.5500 ;
      RECT 0.0000 295.5500 695.6000 299.2500 ;
      RECT 0.7000 295.2500 695.6000 295.5500 ;
      RECT 0.0000 291.5500 695.6000 295.2500 ;
      RECT 0.7000 291.2500 695.6000 291.5500 ;
      RECT 0.0000 287.5500 695.6000 291.2500 ;
      RECT 0.7000 287.2500 695.6000 287.5500 ;
      RECT 0.0000 283.5500 695.6000 287.2500 ;
      RECT 0.7000 283.2500 695.6000 283.5500 ;
      RECT 0.0000 279.5500 695.6000 283.2500 ;
      RECT 0.7000 279.2500 695.6000 279.5500 ;
      RECT 0.0000 275.5500 695.6000 279.2500 ;
      RECT 0.7000 275.2500 695.6000 275.5500 ;
      RECT 0.0000 271.5500 695.6000 275.2500 ;
      RECT 0.7000 271.2500 695.6000 271.5500 ;
      RECT 0.0000 267.5500 695.6000 271.2500 ;
      RECT 0.7000 267.2500 695.6000 267.5500 ;
      RECT 0.0000 263.5500 695.6000 267.2500 ;
      RECT 0.7000 263.2500 695.6000 263.5500 ;
      RECT 0.0000 259.5500 695.6000 263.2500 ;
      RECT 0.7000 259.2500 695.6000 259.5500 ;
      RECT 0.0000 255.5500 695.6000 259.2500 ;
      RECT 0.7000 255.2500 695.6000 255.5500 ;
      RECT 0.0000 251.5500 695.6000 255.2500 ;
      RECT 0.7000 251.2500 695.6000 251.5500 ;
      RECT 0.0000 247.5500 695.6000 251.2500 ;
      RECT 0.7000 247.2500 695.6000 247.5500 ;
      RECT 0.0000 243.5500 695.6000 247.2500 ;
      RECT 0.7000 243.2500 695.6000 243.5500 ;
      RECT 0.0000 239.5500 695.6000 243.2500 ;
      RECT 0.7000 239.2500 695.6000 239.5500 ;
      RECT 0.0000 235.5500 695.6000 239.2500 ;
      RECT 0.7000 235.2500 695.6000 235.5500 ;
      RECT 0.0000 231.5500 695.6000 235.2500 ;
      RECT 0.7000 231.2500 695.6000 231.5500 ;
      RECT 0.0000 227.5500 695.6000 231.2500 ;
      RECT 0.7000 227.2500 695.6000 227.5500 ;
      RECT 0.0000 223.5500 695.6000 227.2500 ;
      RECT 0.7000 223.2500 695.6000 223.5500 ;
      RECT 0.0000 219.5500 695.6000 223.2500 ;
      RECT 0.7000 219.2500 695.6000 219.5500 ;
      RECT 0.0000 215.5500 695.6000 219.2500 ;
      RECT 0.7000 215.2500 695.6000 215.5500 ;
      RECT 0.0000 211.5500 695.6000 215.2500 ;
      RECT 0.7000 211.2500 695.6000 211.5500 ;
      RECT 0.0000 207.5500 695.6000 211.2500 ;
      RECT 0.7000 207.2500 695.6000 207.5500 ;
      RECT 0.0000 203.5500 695.6000 207.2500 ;
      RECT 0.7000 203.2500 695.6000 203.5500 ;
      RECT 0.0000 199.5500 695.6000 203.2500 ;
      RECT 0.7000 199.2500 695.6000 199.5500 ;
      RECT 0.0000 195.5500 695.6000 199.2500 ;
      RECT 0.7000 195.2500 695.6000 195.5500 ;
      RECT 0.0000 191.5500 695.6000 195.2500 ;
      RECT 0.7000 191.2500 695.6000 191.5500 ;
      RECT 0.0000 187.5500 695.6000 191.2500 ;
      RECT 0.7000 187.2500 695.6000 187.5500 ;
      RECT 0.0000 183.5500 695.6000 187.2500 ;
      RECT 0.7000 183.2500 695.6000 183.5500 ;
      RECT 0.0000 179.5500 695.6000 183.2500 ;
      RECT 0.7000 179.2500 695.6000 179.5500 ;
      RECT 0.0000 175.5500 695.6000 179.2500 ;
      RECT 0.7000 175.2500 695.6000 175.5500 ;
      RECT 0.0000 171.5500 695.6000 175.2500 ;
      RECT 0.7000 171.2500 695.6000 171.5500 ;
      RECT 0.0000 167.5500 695.6000 171.2500 ;
      RECT 0.7000 167.2500 695.6000 167.5500 ;
      RECT 0.0000 163.5500 695.6000 167.2500 ;
      RECT 0.7000 163.2500 695.6000 163.5500 ;
      RECT 0.0000 159.5500 695.6000 163.2500 ;
      RECT 0.7000 159.2500 695.6000 159.5500 ;
      RECT 0.0000 155.5500 695.6000 159.2500 ;
      RECT 0.7000 155.2500 695.6000 155.5500 ;
      RECT 0.0000 151.5500 695.6000 155.2500 ;
      RECT 0.7000 151.2500 695.6000 151.5500 ;
      RECT 0.0000 147.5500 695.6000 151.2500 ;
      RECT 0.7000 147.2500 695.6000 147.5500 ;
      RECT 0.0000 143.5500 695.6000 147.2500 ;
      RECT 0.7000 143.2500 695.6000 143.5500 ;
      RECT 0.0000 139.5500 695.6000 143.2500 ;
      RECT 0.7000 139.2500 695.6000 139.5500 ;
      RECT 0.0000 135.5500 695.6000 139.2500 ;
      RECT 0.7000 135.2500 695.6000 135.5500 ;
      RECT 0.0000 131.5500 695.6000 135.2500 ;
      RECT 0.7000 131.2500 695.6000 131.5500 ;
      RECT 0.0000 127.5500 695.6000 131.2500 ;
      RECT 0.7000 127.2500 695.6000 127.5500 ;
      RECT 0.0000 123.5500 695.6000 127.2500 ;
      RECT 0.7000 123.2500 695.6000 123.5500 ;
      RECT 0.0000 119.5500 695.6000 123.2500 ;
      RECT 0.7000 119.2500 695.6000 119.5500 ;
      RECT 0.0000 115.5500 695.6000 119.2500 ;
      RECT 0.7000 115.2500 695.6000 115.5500 ;
      RECT 0.0000 111.5500 695.6000 115.2500 ;
      RECT 0.7000 111.2500 695.6000 111.5500 ;
      RECT 0.0000 107.5500 695.6000 111.2500 ;
      RECT 0.7000 107.2500 695.6000 107.5500 ;
      RECT 0.0000 103.5500 695.6000 107.2500 ;
      RECT 0.7000 103.2500 695.6000 103.5500 ;
      RECT 0.0000 99.5500 695.6000 103.2500 ;
      RECT 0.7000 99.2500 695.6000 99.5500 ;
      RECT 0.0000 95.5500 695.6000 99.2500 ;
      RECT 0.7000 95.2500 695.6000 95.5500 ;
      RECT 0.0000 91.5500 695.6000 95.2500 ;
      RECT 0.7000 91.2500 695.6000 91.5500 ;
      RECT 0.0000 87.5500 695.6000 91.2500 ;
      RECT 0.7000 87.2500 695.6000 87.5500 ;
      RECT 0.0000 83.5500 695.6000 87.2500 ;
      RECT 0.7000 83.2500 695.6000 83.5500 ;
      RECT 0.0000 79.5500 695.6000 83.2500 ;
      RECT 0.7000 79.2500 695.6000 79.5500 ;
      RECT 0.0000 75.5500 695.6000 79.2500 ;
      RECT 0.7000 75.2500 695.6000 75.5500 ;
      RECT 0.0000 71.5500 695.6000 75.2500 ;
      RECT 0.7000 71.2500 695.6000 71.5500 ;
      RECT 0.0000 67.5500 695.6000 71.2500 ;
      RECT 0.7000 67.2500 695.6000 67.5500 ;
      RECT 0.0000 63.5500 695.6000 67.2500 ;
      RECT 0.7000 63.2500 695.6000 63.5500 ;
      RECT 0.0000 59.5500 695.6000 63.2500 ;
      RECT 0.7000 59.2500 695.6000 59.5500 ;
      RECT 0.0000 55.5500 695.6000 59.2500 ;
      RECT 0.7000 55.2500 695.6000 55.5500 ;
      RECT 0.0000 0.0000 695.6000 55.2500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 695.6000 695.0000 ;
  END
END fullchip

END LIBRARY
