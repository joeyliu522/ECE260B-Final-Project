##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Wed Mar 19 04:16:30 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 820.0000 BY 420.0000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 217.7500 0.5200 217.8500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.8500 0.0000 663.9500 0.5200 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.8500 0.0000 659.9500 0.5200 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.8500 0.0000 655.9500 0.5200 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.8500 0.0000 651.9500 0.5200 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.8500 0.0000 647.9500 0.5200 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.8500 0.0000 643.9500 0.5200 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.8500 0.0000 639.9500 0.5200 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.8500 0.0000 635.9500 0.5200 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.8500 0.0000 631.9500 0.5200 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.8500 0.0000 627.9500 0.5200 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.8500 0.0000 623.9500 0.5200 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.8500 0.0000 619.9500 0.5200 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.8500 0.0000 615.9500 0.5200 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.8500 0.0000 611.9500 0.5200 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.8500 0.0000 607.9500 0.5200 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.8500 0.0000 603.9500 0.5200 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.8500 0.0000 599.9500 0.5200 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.8500 0.0000 595.9500 0.5200 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.8500 0.0000 591.9500 0.5200 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.8500 0.0000 587.9500 0.5200 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.8500 0.0000 583.9500 0.5200 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 0.0000 579.9500 0.5200 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.8500 0.0000 575.9500 0.5200 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.8500 0.0000 571.9500 0.5200 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.8500 0.0000 567.9500 0.5200 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.8500 0.0000 563.9500 0.5200 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.8500 0.0000 559.9500 0.5200 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.8500 0.0000 555.9500 0.5200 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.8500 0.0000 551.9500 0.5200 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.8500 0.0000 547.9500 0.5200 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 0.0000 543.9500 0.5200 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.8500 0.0000 539.9500 0.5200 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 0.0000 535.9500 0.5200 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.8500 0.0000 531.9500 0.5200 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.8500 0.0000 527.9500 0.5200 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.8500 0.0000 523.9500 0.5200 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.8500 0.0000 519.9500 0.5200 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.8500 0.0000 515.9500 0.5200 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.8500 0.0000 511.9500 0.5200 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 0.0000 507.9500 0.5200 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.8500 0.0000 503.9500 0.5200 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.8500 0.0000 499.9500 0.5200 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.8500 0.0000 495.9500 0.5200 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.8500 0.0000 491.9500 0.5200 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.8500 0.0000 487.9500 0.5200 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.8500 0.0000 483.9500 0.5200 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.8500 0.0000 479.9500 0.5200 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.8500 0.0000 475.9500 0.5200 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.8500 0.0000 471.9500 0.5200 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.8500 0.0000 467.9500 0.5200 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.8500 0.0000 463.9500 0.5200 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.8500 0.0000 459.9500 0.5200 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.8500 0.0000 455.9500 0.5200 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.8500 0.0000 451.9500 0.5200 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.8500 0.0000 447.9500 0.5200 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.8500 0.0000 443.9500 0.5200 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.8500 0.0000 439.9500 0.5200 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.8500 0.0000 435.9500 0.5200 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.8500 0.0000 431.9500 0.5200 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.8500 0.0000 427.9500 0.5200 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.8500 0.0000 423.9500 0.5200 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.8500 0.0000 419.9500 0.5200 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.8500 0.0000 415.9500 0.5200 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.8500 0.0000 411.9500 0.5200 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.8500 0.0000 407.9500 0.5200 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.8500 0.0000 403.9500 0.5200 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.8500 0.0000 399.9500 0.5200 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.8500 0.0000 395.9500 0.5200 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.8500 0.0000 391.9500 0.5200 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.8500 0.0000 387.9500 0.5200 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.8500 0.0000 383.9500 0.5200 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.8500 0.0000 379.9500 0.5200 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.8500 0.0000 375.9500 0.5200 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.8500 0.0000 371.9500 0.5200 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.8500 0.0000 367.9500 0.5200 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.8500 0.0000 363.9500 0.5200 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.8500 0.0000 359.9500 0.5200 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.8500 0.0000 355.9500 0.5200 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.8500 0.0000 351.9500 0.5200 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.8500 0.0000 347.9500 0.5200 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.8500 0.0000 343.9500 0.5200 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.8500 0.0000 339.9500 0.5200 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.8500 0.0000 335.9500 0.5200 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.8500 0.0000 331.9500 0.5200 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.8500 0.0000 327.9500 0.5200 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.8500 0.0000 323.9500 0.5200 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.8500 0.0000 319.9500 0.5200 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.8500 0.0000 315.9500 0.5200 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.8500 0.0000 311.9500 0.5200 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.8500 0.0000 307.9500 0.5200 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.8500 0.0000 303.9500 0.5200 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.8500 0.0000 299.9500 0.5200 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.8500 0.0000 295.9500 0.5200 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.8500 0.0000 291.9500 0.5200 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.8500 0.0000 287.9500 0.5200 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.8500 0.0000 283.9500 0.5200 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.8500 0.0000 279.9500 0.5200 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.8500 0.0000 275.9500 0.5200 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.8500 0.0000 271.9500 0.5200 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.8500 0.0000 267.9500 0.5200 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.8500 0.0000 263.9500 0.5200 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.8500 0.0000 259.9500 0.5200 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.8500 0.0000 255.9500 0.5200 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.8500 0.0000 251.9500 0.5200 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.8500 0.0000 247.9500 0.5200 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.8500 0.0000 243.9500 0.5200 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.8500 0.0000 239.9500 0.5200 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.8500 0.0000 235.9500 0.5200 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.8500 0.0000 231.9500 0.5200 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.8500 0.0000 227.9500 0.5200 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.8500 0.0000 223.9500 0.5200 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.8500 0.0000 219.9500 0.5200 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.8500 0.0000 215.9500 0.5200 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.8500 0.0000 211.9500 0.5200 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.8500 0.0000 207.9500 0.5200 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.8500 0.0000 203.9500 0.5200 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.8500 0.0000 199.9500 0.5200 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.8500 0.0000 195.9500 0.5200 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.8500 0.0000 191.9500 0.5200 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.8500 0.0000 187.9500 0.5200 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.8500 0.0000 183.9500 0.5200 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.8500 0.0000 179.9500 0.5200 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.8500 0.0000 175.9500 0.5200 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.8500 0.0000 171.9500 0.5200 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.8500 0.0000 167.9500 0.5200 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 0.0000 163.9500 0.5200 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.8500 0.0000 159.9500 0.5200 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 0.0000 155.9500 0.5200 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.8500 419.4800 663.9500 420.0000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.8500 419.4800 659.9500 420.0000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.8500 419.4800 655.9500 420.0000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.8500 419.4800 651.9500 420.0000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.8500 419.4800 647.9500 420.0000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.8500 419.4800 643.9500 420.0000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.8500 419.4800 639.9500 420.0000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.8500 419.4800 635.9500 420.0000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.8500 419.4800 631.9500 420.0000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.8500 419.4800 627.9500 420.0000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.8500 419.4800 623.9500 420.0000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.8500 419.4800 619.9500 420.0000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.8500 419.4800 615.9500 420.0000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.8500 419.4800 611.9500 420.0000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.8500 419.4800 607.9500 420.0000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.8500 419.4800 603.9500 420.0000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.8500 419.4800 599.9500 420.0000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.8500 419.4800 595.9500 420.0000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.8500 419.4800 591.9500 420.0000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.8500 419.4800 587.9500 420.0000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.8500 419.4800 583.9500 420.0000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 419.4800 579.9500 420.0000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.8500 419.4800 575.9500 420.0000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.8500 419.4800 571.9500 420.0000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.8500 419.4800 567.9500 420.0000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.8500 419.4800 563.9500 420.0000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.8500 419.4800 559.9500 420.0000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.8500 419.4800 555.9500 420.0000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.8500 419.4800 551.9500 420.0000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.8500 419.4800 547.9500 420.0000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 419.4800 543.9500 420.0000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.8500 419.4800 539.9500 420.0000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 419.4800 535.9500 420.0000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.8500 419.4800 531.9500 420.0000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.8500 419.4800 527.9500 420.0000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.8500 419.4800 523.9500 420.0000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.8500 419.4800 519.9500 420.0000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.8500 419.4800 515.9500 420.0000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.8500 419.4800 511.9500 420.0000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 419.4800 507.9500 420.0000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.8500 419.4800 503.9500 420.0000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.8500 419.4800 499.9500 420.0000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.8500 419.4800 495.9500 420.0000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.8500 419.4800 491.9500 420.0000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.8500 419.4800 487.9500 420.0000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.8500 419.4800 483.9500 420.0000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.8500 419.4800 479.9500 420.0000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.8500 419.4800 475.9500 420.0000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.8500 419.4800 471.9500 420.0000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.8500 419.4800 467.9500 420.0000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.8500 419.4800 463.9500 420.0000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.8500 419.4800 459.9500 420.0000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.8500 419.4800 455.9500 420.0000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.8500 419.4800 451.9500 420.0000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.8500 419.4800 447.9500 420.0000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.8500 419.4800 443.9500 420.0000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.8500 419.4800 439.9500 420.0000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.8500 419.4800 435.9500 420.0000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.8500 419.4800 431.9500 420.0000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.8500 419.4800 427.9500 420.0000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.8500 419.4800 423.9500 420.0000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.8500 419.4800 419.9500 420.0000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.8500 419.4800 415.9500 420.0000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.8500 419.4800 411.9500 420.0000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.8500 419.4800 407.9500 420.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.8500 419.4800 403.9500 420.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.8500 419.4800 399.9500 420.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.8500 419.4800 395.9500 420.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.8500 419.4800 391.9500 420.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.8500 419.4800 387.9500 420.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.8500 419.4800 383.9500 420.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.8500 419.4800 379.9500 420.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.8500 419.4800 375.9500 420.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.8500 419.4800 371.9500 420.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.8500 419.4800 367.9500 420.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.8500 419.4800 363.9500 420.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.8500 419.4800 359.9500 420.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.8500 419.4800 355.9500 420.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.8500 419.4800 351.9500 420.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.8500 419.4800 347.9500 420.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.8500 419.4800 343.9500 420.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.8500 419.4800 339.9500 420.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.8500 419.4800 335.9500 420.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.8500 419.4800 331.9500 420.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.8500 419.4800 327.9500 420.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.8500 419.4800 323.9500 420.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.8500 419.4800 319.9500 420.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.8500 419.4800 315.9500 420.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.8500 419.4800 311.9500 420.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.8500 419.4800 307.9500 420.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.8500 419.4800 303.9500 420.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.8500 419.4800 299.9500 420.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.8500 419.4800 295.9500 420.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.8500 419.4800 291.9500 420.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.8500 419.4800 287.9500 420.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.8500 419.4800 283.9500 420.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.8500 419.4800 279.9500 420.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.8500 419.4800 275.9500 420.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.8500 419.4800 271.9500 420.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.8500 419.4800 267.9500 420.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.8500 419.4800 263.9500 420.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.8500 419.4800 259.9500 420.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.8500 419.4800 255.9500 420.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.8500 419.4800 251.9500 420.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.8500 419.4800 247.9500 420.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.8500 419.4800 243.9500 420.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.8500 419.4800 239.9500 420.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.8500 419.4800 235.9500 420.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.8500 419.4800 231.9500 420.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.8500 419.4800 227.9500 420.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.8500 419.4800 223.9500 420.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.8500 419.4800 219.9500 420.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.8500 419.4800 215.9500 420.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.8500 419.4800 211.9500 420.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.8500 419.4800 207.9500 420.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.8500 419.4800 203.9500 420.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.8500 419.4800 199.9500 420.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.8500 419.4800 195.9500 420.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.8500 419.4800 191.9500 420.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.8500 419.4800 187.9500 420.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.8500 419.4800 183.9500 420.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.8500 419.4800 179.9500 420.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.8500 419.4800 175.9500 420.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.8500 419.4800 171.9500 420.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.8500 419.4800 167.9500 420.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 419.4800 163.9500 420.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.8500 419.4800 159.9500 420.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 419.4800 155.9500 420.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.7500 0.5200 213.8500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 221.7500 0.5200 221.8500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.7500 0.5200 209.8500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.7500 0.5200 205.8500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.7500 0.5200 201.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 197.7500 0.5200 197.8500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 806.9850 10.0000 807.9850 410.0000 ;
        RECT 693.1300 10.0000 694.1300 410.0000 ;
        RECT 579.2750 10.0000 580.2750 410.0000 ;
        RECT 465.4200 10.0000 466.4200 410.0000 ;
        RECT 351.5650 10.0000 352.5650 410.0000 ;
        RECT 237.7100 10.0000 238.7100 410.0000 ;
        RECT 123.8550 10.0000 124.8550 410.0000 ;
        RECT 10.0000 10.0000 11.0000 410.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 808.9850 10.0000 809.9850 410.0000 ;
        RECT 695.1300 10.0000 696.1300 410.0000 ;
        RECT 581.2750 10.0000 582.2750 410.0000 ;
        RECT 467.4200 10.0000 468.4200 410.0000 ;
        RECT 353.5650 10.0000 354.5650 410.0000 ;
        RECT 239.7100 10.0000 240.7100 410.0000 ;
        RECT 125.8550 10.0000 126.8550 410.0000 ;
        RECT 12.0000 10.0000 13.0000 410.0000 ;
        RECT 12.0000 9.8350 13.0000 10.1650 ;
        RECT 125.8550 9.8350 126.8550 10.1650 ;
        RECT 239.7100 9.8350 240.7100 10.1650 ;
        RECT 353.5650 9.8350 354.5650 10.1650 ;
        RECT 467.4200 9.8350 468.4200 10.1650 ;
        RECT 581.2750 9.8350 582.2750 10.1650 ;
        RECT 695.1300 9.8350 696.1300 10.1650 ;
        RECT 808.9850 9.8350 809.9850 10.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 820.0000 420.0000 ;
    LAYER M2 ;
      RECT 664.0500 419.3800 820.0000 420.0000 ;
      RECT 660.0500 419.3800 663.7500 420.0000 ;
      RECT 656.0500 419.3800 659.7500 420.0000 ;
      RECT 652.0500 419.3800 655.7500 420.0000 ;
      RECT 648.0500 419.3800 651.7500 420.0000 ;
      RECT 644.0500 419.3800 647.7500 420.0000 ;
      RECT 640.0500 419.3800 643.7500 420.0000 ;
      RECT 636.0500 419.3800 639.7500 420.0000 ;
      RECT 632.0500 419.3800 635.7500 420.0000 ;
      RECT 628.0500 419.3800 631.7500 420.0000 ;
      RECT 624.0500 419.3800 627.7500 420.0000 ;
      RECT 620.0500 419.3800 623.7500 420.0000 ;
      RECT 616.0500 419.3800 619.7500 420.0000 ;
      RECT 612.0500 419.3800 615.7500 420.0000 ;
      RECT 608.0500 419.3800 611.7500 420.0000 ;
      RECT 604.0500 419.3800 607.7500 420.0000 ;
      RECT 600.0500 419.3800 603.7500 420.0000 ;
      RECT 596.0500 419.3800 599.7500 420.0000 ;
      RECT 592.0500 419.3800 595.7500 420.0000 ;
      RECT 588.0500 419.3800 591.7500 420.0000 ;
      RECT 584.0500 419.3800 587.7500 420.0000 ;
      RECT 580.0500 419.3800 583.7500 420.0000 ;
      RECT 576.0500 419.3800 579.7500 420.0000 ;
      RECT 572.0500 419.3800 575.7500 420.0000 ;
      RECT 568.0500 419.3800 571.7500 420.0000 ;
      RECT 564.0500 419.3800 567.7500 420.0000 ;
      RECT 560.0500 419.3800 563.7500 420.0000 ;
      RECT 556.0500 419.3800 559.7500 420.0000 ;
      RECT 552.0500 419.3800 555.7500 420.0000 ;
      RECT 548.0500 419.3800 551.7500 420.0000 ;
      RECT 544.0500 419.3800 547.7500 420.0000 ;
      RECT 540.0500 419.3800 543.7500 420.0000 ;
      RECT 536.0500 419.3800 539.7500 420.0000 ;
      RECT 532.0500 419.3800 535.7500 420.0000 ;
      RECT 528.0500 419.3800 531.7500 420.0000 ;
      RECT 524.0500 419.3800 527.7500 420.0000 ;
      RECT 520.0500 419.3800 523.7500 420.0000 ;
      RECT 516.0500 419.3800 519.7500 420.0000 ;
      RECT 512.0500 419.3800 515.7500 420.0000 ;
      RECT 508.0500 419.3800 511.7500 420.0000 ;
      RECT 504.0500 419.3800 507.7500 420.0000 ;
      RECT 500.0500 419.3800 503.7500 420.0000 ;
      RECT 496.0500 419.3800 499.7500 420.0000 ;
      RECT 492.0500 419.3800 495.7500 420.0000 ;
      RECT 488.0500 419.3800 491.7500 420.0000 ;
      RECT 484.0500 419.3800 487.7500 420.0000 ;
      RECT 480.0500 419.3800 483.7500 420.0000 ;
      RECT 476.0500 419.3800 479.7500 420.0000 ;
      RECT 472.0500 419.3800 475.7500 420.0000 ;
      RECT 468.0500 419.3800 471.7500 420.0000 ;
      RECT 464.0500 419.3800 467.7500 420.0000 ;
      RECT 460.0500 419.3800 463.7500 420.0000 ;
      RECT 456.0500 419.3800 459.7500 420.0000 ;
      RECT 452.0500 419.3800 455.7500 420.0000 ;
      RECT 448.0500 419.3800 451.7500 420.0000 ;
      RECT 444.0500 419.3800 447.7500 420.0000 ;
      RECT 440.0500 419.3800 443.7500 420.0000 ;
      RECT 436.0500 419.3800 439.7500 420.0000 ;
      RECT 432.0500 419.3800 435.7500 420.0000 ;
      RECT 428.0500 419.3800 431.7500 420.0000 ;
      RECT 424.0500 419.3800 427.7500 420.0000 ;
      RECT 420.0500 419.3800 423.7500 420.0000 ;
      RECT 416.0500 419.3800 419.7500 420.0000 ;
      RECT 412.0500 419.3800 415.7500 420.0000 ;
      RECT 408.0500 419.3800 411.7500 420.0000 ;
      RECT 404.0500 419.3800 407.7500 420.0000 ;
      RECT 400.0500 419.3800 403.7500 420.0000 ;
      RECT 396.0500 419.3800 399.7500 420.0000 ;
      RECT 392.0500 419.3800 395.7500 420.0000 ;
      RECT 388.0500 419.3800 391.7500 420.0000 ;
      RECT 384.0500 419.3800 387.7500 420.0000 ;
      RECT 380.0500 419.3800 383.7500 420.0000 ;
      RECT 376.0500 419.3800 379.7500 420.0000 ;
      RECT 372.0500 419.3800 375.7500 420.0000 ;
      RECT 368.0500 419.3800 371.7500 420.0000 ;
      RECT 364.0500 419.3800 367.7500 420.0000 ;
      RECT 360.0500 419.3800 363.7500 420.0000 ;
      RECT 356.0500 419.3800 359.7500 420.0000 ;
      RECT 352.0500 419.3800 355.7500 420.0000 ;
      RECT 348.0500 419.3800 351.7500 420.0000 ;
      RECT 344.0500 419.3800 347.7500 420.0000 ;
      RECT 340.0500 419.3800 343.7500 420.0000 ;
      RECT 336.0500 419.3800 339.7500 420.0000 ;
      RECT 332.0500 419.3800 335.7500 420.0000 ;
      RECT 328.0500 419.3800 331.7500 420.0000 ;
      RECT 324.0500 419.3800 327.7500 420.0000 ;
      RECT 320.0500 419.3800 323.7500 420.0000 ;
      RECT 316.0500 419.3800 319.7500 420.0000 ;
      RECT 312.0500 419.3800 315.7500 420.0000 ;
      RECT 308.0500 419.3800 311.7500 420.0000 ;
      RECT 304.0500 419.3800 307.7500 420.0000 ;
      RECT 300.0500 419.3800 303.7500 420.0000 ;
      RECT 296.0500 419.3800 299.7500 420.0000 ;
      RECT 292.0500 419.3800 295.7500 420.0000 ;
      RECT 288.0500 419.3800 291.7500 420.0000 ;
      RECT 284.0500 419.3800 287.7500 420.0000 ;
      RECT 280.0500 419.3800 283.7500 420.0000 ;
      RECT 276.0500 419.3800 279.7500 420.0000 ;
      RECT 272.0500 419.3800 275.7500 420.0000 ;
      RECT 268.0500 419.3800 271.7500 420.0000 ;
      RECT 264.0500 419.3800 267.7500 420.0000 ;
      RECT 260.0500 419.3800 263.7500 420.0000 ;
      RECT 256.0500 419.3800 259.7500 420.0000 ;
      RECT 252.0500 419.3800 255.7500 420.0000 ;
      RECT 248.0500 419.3800 251.7500 420.0000 ;
      RECT 244.0500 419.3800 247.7500 420.0000 ;
      RECT 240.0500 419.3800 243.7500 420.0000 ;
      RECT 236.0500 419.3800 239.7500 420.0000 ;
      RECT 232.0500 419.3800 235.7500 420.0000 ;
      RECT 228.0500 419.3800 231.7500 420.0000 ;
      RECT 224.0500 419.3800 227.7500 420.0000 ;
      RECT 220.0500 419.3800 223.7500 420.0000 ;
      RECT 216.0500 419.3800 219.7500 420.0000 ;
      RECT 212.0500 419.3800 215.7500 420.0000 ;
      RECT 208.0500 419.3800 211.7500 420.0000 ;
      RECT 204.0500 419.3800 207.7500 420.0000 ;
      RECT 200.0500 419.3800 203.7500 420.0000 ;
      RECT 196.0500 419.3800 199.7500 420.0000 ;
      RECT 192.0500 419.3800 195.7500 420.0000 ;
      RECT 188.0500 419.3800 191.7500 420.0000 ;
      RECT 184.0500 419.3800 187.7500 420.0000 ;
      RECT 180.0500 419.3800 183.7500 420.0000 ;
      RECT 176.0500 419.3800 179.7500 420.0000 ;
      RECT 172.0500 419.3800 175.7500 420.0000 ;
      RECT 168.0500 419.3800 171.7500 420.0000 ;
      RECT 164.0500 419.3800 167.7500 420.0000 ;
      RECT 160.0500 419.3800 163.7500 420.0000 ;
      RECT 156.0500 419.3800 159.7500 420.0000 ;
      RECT 0.0000 419.3800 155.7500 420.0000 ;
      RECT 0.0000 0.6200 820.0000 419.3800 ;
      RECT 664.0500 0.0000 820.0000 0.6200 ;
      RECT 660.0500 0.0000 663.7500 0.6200 ;
      RECT 656.0500 0.0000 659.7500 0.6200 ;
      RECT 652.0500 0.0000 655.7500 0.6200 ;
      RECT 648.0500 0.0000 651.7500 0.6200 ;
      RECT 644.0500 0.0000 647.7500 0.6200 ;
      RECT 640.0500 0.0000 643.7500 0.6200 ;
      RECT 636.0500 0.0000 639.7500 0.6200 ;
      RECT 632.0500 0.0000 635.7500 0.6200 ;
      RECT 628.0500 0.0000 631.7500 0.6200 ;
      RECT 624.0500 0.0000 627.7500 0.6200 ;
      RECT 620.0500 0.0000 623.7500 0.6200 ;
      RECT 616.0500 0.0000 619.7500 0.6200 ;
      RECT 612.0500 0.0000 615.7500 0.6200 ;
      RECT 608.0500 0.0000 611.7500 0.6200 ;
      RECT 604.0500 0.0000 607.7500 0.6200 ;
      RECT 600.0500 0.0000 603.7500 0.6200 ;
      RECT 596.0500 0.0000 599.7500 0.6200 ;
      RECT 592.0500 0.0000 595.7500 0.6200 ;
      RECT 588.0500 0.0000 591.7500 0.6200 ;
      RECT 584.0500 0.0000 587.7500 0.6200 ;
      RECT 580.0500 0.0000 583.7500 0.6200 ;
      RECT 576.0500 0.0000 579.7500 0.6200 ;
      RECT 572.0500 0.0000 575.7500 0.6200 ;
      RECT 568.0500 0.0000 571.7500 0.6200 ;
      RECT 564.0500 0.0000 567.7500 0.6200 ;
      RECT 560.0500 0.0000 563.7500 0.6200 ;
      RECT 556.0500 0.0000 559.7500 0.6200 ;
      RECT 552.0500 0.0000 555.7500 0.6200 ;
      RECT 548.0500 0.0000 551.7500 0.6200 ;
      RECT 544.0500 0.0000 547.7500 0.6200 ;
      RECT 540.0500 0.0000 543.7500 0.6200 ;
      RECT 536.0500 0.0000 539.7500 0.6200 ;
      RECT 532.0500 0.0000 535.7500 0.6200 ;
      RECT 528.0500 0.0000 531.7500 0.6200 ;
      RECT 524.0500 0.0000 527.7500 0.6200 ;
      RECT 520.0500 0.0000 523.7500 0.6200 ;
      RECT 516.0500 0.0000 519.7500 0.6200 ;
      RECT 512.0500 0.0000 515.7500 0.6200 ;
      RECT 508.0500 0.0000 511.7500 0.6200 ;
      RECT 504.0500 0.0000 507.7500 0.6200 ;
      RECT 500.0500 0.0000 503.7500 0.6200 ;
      RECT 496.0500 0.0000 499.7500 0.6200 ;
      RECT 492.0500 0.0000 495.7500 0.6200 ;
      RECT 488.0500 0.0000 491.7500 0.6200 ;
      RECT 484.0500 0.0000 487.7500 0.6200 ;
      RECT 480.0500 0.0000 483.7500 0.6200 ;
      RECT 476.0500 0.0000 479.7500 0.6200 ;
      RECT 472.0500 0.0000 475.7500 0.6200 ;
      RECT 468.0500 0.0000 471.7500 0.6200 ;
      RECT 464.0500 0.0000 467.7500 0.6200 ;
      RECT 460.0500 0.0000 463.7500 0.6200 ;
      RECT 456.0500 0.0000 459.7500 0.6200 ;
      RECT 452.0500 0.0000 455.7500 0.6200 ;
      RECT 448.0500 0.0000 451.7500 0.6200 ;
      RECT 444.0500 0.0000 447.7500 0.6200 ;
      RECT 440.0500 0.0000 443.7500 0.6200 ;
      RECT 436.0500 0.0000 439.7500 0.6200 ;
      RECT 432.0500 0.0000 435.7500 0.6200 ;
      RECT 428.0500 0.0000 431.7500 0.6200 ;
      RECT 424.0500 0.0000 427.7500 0.6200 ;
      RECT 420.0500 0.0000 423.7500 0.6200 ;
      RECT 416.0500 0.0000 419.7500 0.6200 ;
      RECT 412.0500 0.0000 415.7500 0.6200 ;
      RECT 408.0500 0.0000 411.7500 0.6200 ;
      RECT 404.0500 0.0000 407.7500 0.6200 ;
      RECT 400.0500 0.0000 403.7500 0.6200 ;
      RECT 396.0500 0.0000 399.7500 0.6200 ;
      RECT 392.0500 0.0000 395.7500 0.6200 ;
      RECT 388.0500 0.0000 391.7500 0.6200 ;
      RECT 384.0500 0.0000 387.7500 0.6200 ;
      RECT 380.0500 0.0000 383.7500 0.6200 ;
      RECT 376.0500 0.0000 379.7500 0.6200 ;
      RECT 372.0500 0.0000 375.7500 0.6200 ;
      RECT 368.0500 0.0000 371.7500 0.6200 ;
      RECT 364.0500 0.0000 367.7500 0.6200 ;
      RECT 360.0500 0.0000 363.7500 0.6200 ;
      RECT 356.0500 0.0000 359.7500 0.6200 ;
      RECT 352.0500 0.0000 355.7500 0.6200 ;
      RECT 348.0500 0.0000 351.7500 0.6200 ;
      RECT 344.0500 0.0000 347.7500 0.6200 ;
      RECT 340.0500 0.0000 343.7500 0.6200 ;
      RECT 336.0500 0.0000 339.7500 0.6200 ;
      RECT 332.0500 0.0000 335.7500 0.6200 ;
      RECT 328.0500 0.0000 331.7500 0.6200 ;
      RECT 324.0500 0.0000 327.7500 0.6200 ;
      RECT 320.0500 0.0000 323.7500 0.6200 ;
      RECT 316.0500 0.0000 319.7500 0.6200 ;
      RECT 312.0500 0.0000 315.7500 0.6200 ;
      RECT 308.0500 0.0000 311.7500 0.6200 ;
      RECT 304.0500 0.0000 307.7500 0.6200 ;
      RECT 300.0500 0.0000 303.7500 0.6200 ;
      RECT 296.0500 0.0000 299.7500 0.6200 ;
      RECT 292.0500 0.0000 295.7500 0.6200 ;
      RECT 288.0500 0.0000 291.7500 0.6200 ;
      RECT 284.0500 0.0000 287.7500 0.6200 ;
      RECT 280.0500 0.0000 283.7500 0.6200 ;
      RECT 276.0500 0.0000 279.7500 0.6200 ;
      RECT 272.0500 0.0000 275.7500 0.6200 ;
      RECT 268.0500 0.0000 271.7500 0.6200 ;
      RECT 264.0500 0.0000 267.7500 0.6200 ;
      RECT 260.0500 0.0000 263.7500 0.6200 ;
      RECT 256.0500 0.0000 259.7500 0.6200 ;
      RECT 252.0500 0.0000 255.7500 0.6200 ;
      RECT 248.0500 0.0000 251.7500 0.6200 ;
      RECT 244.0500 0.0000 247.7500 0.6200 ;
      RECT 240.0500 0.0000 243.7500 0.6200 ;
      RECT 236.0500 0.0000 239.7500 0.6200 ;
      RECT 232.0500 0.0000 235.7500 0.6200 ;
      RECT 228.0500 0.0000 231.7500 0.6200 ;
      RECT 224.0500 0.0000 227.7500 0.6200 ;
      RECT 220.0500 0.0000 223.7500 0.6200 ;
      RECT 216.0500 0.0000 219.7500 0.6200 ;
      RECT 212.0500 0.0000 215.7500 0.6200 ;
      RECT 208.0500 0.0000 211.7500 0.6200 ;
      RECT 204.0500 0.0000 207.7500 0.6200 ;
      RECT 200.0500 0.0000 203.7500 0.6200 ;
      RECT 196.0500 0.0000 199.7500 0.6200 ;
      RECT 192.0500 0.0000 195.7500 0.6200 ;
      RECT 188.0500 0.0000 191.7500 0.6200 ;
      RECT 184.0500 0.0000 187.7500 0.6200 ;
      RECT 180.0500 0.0000 183.7500 0.6200 ;
      RECT 176.0500 0.0000 179.7500 0.6200 ;
      RECT 172.0500 0.0000 175.7500 0.6200 ;
      RECT 168.0500 0.0000 171.7500 0.6200 ;
      RECT 164.0500 0.0000 167.7500 0.6200 ;
      RECT 160.0500 0.0000 163.7500 0.6200 ;
      RECT 156.0500 0.0000 159.7500 0.6200 ;
      RECT 0.0000 0.0000 155.7500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 221.9500 820.0000 420.0000 ;
      RECT 0.6200 221.6500 820.0000 221.9500 ;
      RECT 0.0000 217.9500 820.0000 221.6500 ;
      RECT 0.6200 217.6500 820.0000 217.9500 ;
      RECT 0.0000 213.9500 820.0000 217.6500 ;
      RECT 0.6200 213.6500 820.0000 213.9500 ;
      RECT 0.0000 209.9500 820.0000 213.6500 ;
      RECT 0.6200 209.6500 820.0000 209.9500 ;
      RECT 0.0000 205.9500 820.0000 209.6500 ;
      RECT 0.6200 205.6500 820.0000 205.9500 ;
      RECT 0.0000 201.9500 820.0000 205.6500 ;
      RECT 0.6200 201.6500 820.0000 201.9500 ;
      RECT 0.0000 197.9500 820.0000 201.6500 ;
      RECT 0.6200 197.6500 820.0000 197.9500 ;
      RECT 0.0000 0.0000 820.0000 197.6500 ;
    LAYER M4 ;
      RECT 0.0000 410.1600 820.0000 420.0000 ;
      RECT 808.1450 9.8400 808.8250 410.1600 ;
      RECT 696.2900 9.8400 806.8250 410.1600 ;
      RECT 694.2900 9.8400 694.9700 410.1600 ;
      RECT 582.4350 9.8400 692.9700 410.1600 ;
      RECT 580.4350 9.8400 581.1150 410.1600 ;
      RECT 468.5800 9.8400 579.1150 410.1600 ;
      RECT 466.5800 9.8400 467.2600 410.1600 ;
      RECT 354.7250 9.8400 465.2600 410.1600 ;
      RECT 352.7250 9.8400 353.4050 410.1600 ;
      RECT 240.8700 9.8400 351.4050 410.1600 ;
      RECT 238.8700 9.8400 239.5500 410.1600 ;
      RECT 127.0150 9.8400 237.5500 410.1600 ;
      RECT 125.0150 9.8400 125.6950 410.1600 ;
      RECT 13.1600 9.8400 123.6950 410.1600 ;
      RECT 11.1600 9.8400 11.8400 410.1600 ;
      RECT 0.0000 9.8400 9.8400 410.1600 ;
      RECT 810.1450 9.6750 820.0000 410.1600 ;
      RECT 696.2900 9.6750 808.8250 9.8400 ;
      RECT 582.4350 9.6750 694.9700 9.8400 ;
      RECT 468.5800 9.6750 581.1150 9.8400 ;
      RECT 354.7250 9.6750 467.2600 9.8400 ;
      RECT 240.8700 9.6750 353.4050 9.8400 ;
      RECT 127.0150 9.6750 239.5500 9.8400 ;
      RECT 13.1600 9.6750 125.6950 9.8400 ;
      RECT 0.0000 9.6750 11.8400 9.8400 ;
      RECT 0.0000 0.0000 820.0000 9.6750 ;
  END
END sram_w16

END LIBRARY
