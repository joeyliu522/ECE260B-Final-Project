/home/linux/ieng6/oce/0m/maquilina/Desktop/ece260b/project/Part4/pnr_core/subckt/sram_w16.lef