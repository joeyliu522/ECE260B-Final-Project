##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 14:40:16 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1420.0000 BY 1620.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 809.7500 0.5200 809.8500 ;
    END
  END clk
  PIN sum_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1155.7500 0.5200 1155.8500 ;
    END
  END sum_in[23]
  PIN sum_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1151.7500 0.5200 1151.8500 ;
    END
  END sum_in[22]
  PIN sum_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1147.7500 0.5200 1147.8500 ;
    END
  END sum_in[21]
  PIN sum_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1143.7500 0.5200 1143.8500 ;
    END
  END sum_in[20]
  PIN sum_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1139.7500 0.5200 1139.8500 ;
    END
  END sum_in[19]
  PIN sum_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1135.7500 0.5200 1135.8500 ;
    END
  END sum_in[18]
  PIN sum_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1131.7500 0.5200 1131.8500 ;
    END
  END sum_in[17]
  PIN sum_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1127.7500 0.5200 1127.8500 ;
    END
  END sum_in[16]
  PIN sum_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1123.7500 0.5200 1123.8500 ;
    END
  END sum_in[15]
  PIN sum_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1119.7500 0.5200 1119.8500 ;
    END
  END sum_in[14]
  PIN sum_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1115.7500 0.5200 1115.8500 ;
    END
  END sum_in[13]
  PIN sum_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1111.7500 0.5200 1111.8500 ;
    END
  END sum_in[12]
  PIN sum_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1107.7500 0.5200 1107.8500 ;
    END
  END sum_in[11]
  PIN sum_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1103.7500 0.5200 1103.8500 ;
    END
  END sum_in[10]
  PIN sum_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1099.7500 0.5200 1099.8500 ;
    END
  END sum_in[9]
  PIN sum_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1095.7500 0.5200 1095.8500 ;
    END
  END sum_in[8]
  PIN sum_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1091.7500 0.5200 1091.8500 ;
    END
  END sum_in[7]
  PIN sum_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1087.7500 0.5200 1087.8500 ;
    END
  END sum_in[6]
  PIN sum_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1083.7500 0.5200 1083.8500 ;
    END
  END sum_in[5]
  PIN sum_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1079.7500 0.5200 1079.8500 ;
    END
  END sum_in[4]
  PIN sum_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1075.7500 0.5200 1075.8500 ;
    END
  END sum_in[3]
  PIN sum_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1071.7500 0.5200 1071.8500 ;
    END
  END sum_in[2]
  PIN sum_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1067.7500 0.5200 1067.8500 ;
    END
  END sum_in[1]
  PIN sum_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1063.7500 0.5200 1063.8500 ;
    END
  END sum_in[0]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 764.1500 1420.0000 764.2500 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 768.1500 1420.0000 768.2500 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 772.1500 1420.0000 772.2500 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 776.1500 1420.0000 776.2500 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 780.1500 1420.0000 780.2500 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 784.1500 1420.0000 784.2500 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 788.1500 1420.0000 788.2500 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 792.1500 1420.0000 792.2500 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 796.1500 1420.0000 796.2500 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 800.1500 1420.0000 800.2500 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 804.1500 1420.0000 804.2500 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 808.1500 1420.0000 808.2500 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 812.1500 1420.0000 812.2500 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 816.1500 1420.0000 816.2500 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 820.1500 1420.0000 820.2500 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 824.1500 1420.0000 824.2500 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 828.1500 1420.0000 828.2500 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 832.1500 1420.0000 832.2500 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 836.1500 1420.0000 836.2500 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 840.1500 1420.0000 840.2500 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 844.1500 1420.0000 844.2500 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 848.1500 1420.0000 848.2500 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 852.1500 1420.0000 852.2500 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 856.1500 1420.0000 856.2500 ;
    END
  END sum_out[0]
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 979.7500 0.5200 979.8500 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 975.7500 0.5200 975.8500 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 971.7500 0.5200 971.8500 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 967.7500 0.5200 967.8500 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 963.7500 0.5200 963.8500 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 959.7500 0.5200 959.8500 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 955.7500 0.5200 955.8500 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 951.7500 0.5200 951.8500 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 947.7500 0.5200 947.8500 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 943.7500 0.5200 943.8500 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 939.7500 0.5200 939.8500 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 935.7500 0.5200 935.8500 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 931.7500 0.5200 931.8500 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 927.7500 0.5200 927.8500 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 923.7500 0.5200 923.8500 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 919.7500 0.5200 919.8500 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 915.7500 0.5200 915.8500 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 911.7500 0.5200 911.8500 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 907.7500 0.5200 907.8500 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 903.7500 0.5200 903.8500 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 899.7500 0.5200 899.8500 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 895.7500 0.5200 895.8500 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 891.7500 0.5200 891.8500 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 887.7500 0.5200 887.8500 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 883.7500 0.5200 883.8500 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 879.7500 0.5200 879.8500 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 875.7500 0.5200 875.8500 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 871.7500 0.5200 871.8500 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 867.7500 0.5200 867.8500 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 863.7500 0.5200 863.8500 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 859.7500 0.5200 859.8500 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 855.7500 0.5200 855.8500 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 851.7500 0.5200 851.8500 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 847.7500 0.5200 847.8500 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 843.7500 0.5200 843.8500 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 839.7500 0.5200 839.8500 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 835.7500 0.5200 835.8500 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 831.7500 0.5200 831.8500 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 827.7500 0.5200 827.8500 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 823.7500 0.5200 823.8500 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 819.7500 0.5200 819.8500 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 815.7500 0.5200 815.8500 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 811.7500 0.5200 811.8500 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 807.7500 0.5200 807.8500 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 803.7500 0.5200 803.8500 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 799.7500 0.5200 799.8500 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 795.7500 0.5200 795.8500 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 791.7500 0.5200 791.8500 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 787.7500 0.5200 787.8500 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 783.7500 0.5200 783.8500 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 779.7500 0.5200 779.8500 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 775.7500 0.5200 775.8500 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 771.7500 0.5200 771.8500 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 767.7500 0.5200 767.8500 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 763.7500 0.5200 763.8500 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 759.7500 0.5200 759.8500 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 755.7500 0.5200 755.8500 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 751.7500 0.5200 751.8500 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 747.7500 0.5200 747.8500 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 743.7500 0.5200 743.8500 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 739.7500 0.5200 739.8500 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 735.7500 0.5200 735.8500 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 731.7500 0.5200 731.8500 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 727.7500 0.5200 727.8500 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 723.7500 0.5200 723.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 719.7500 0.5200 719.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 715.7500 0.5200 715.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 711.7500 0.5200 711.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 707.7500 0.5200 707.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 703.7500 0.5200 703.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 699.7500 0.5200 699.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 695.7500 0.5200 695.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 691.7500 0.5200 691.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 687.7500 0.5200 687.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 683.7500 0.5200 683.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 679.7500 0.5200 679.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 675.7500 0.5200 675.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 671.7500 0.5200 671.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 667.7500 0.5200 667.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 663.7500 0.5200 663.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 659.7500 0.5200 659.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 655.7500 0.5200 655.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 651.7500 0.5200 651.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 647.7500 0.5200 647.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 643.7500 0.5200 643.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 639.7500 0.5200 639.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 635.7500 0.5200 635.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 631.7500 0.5200 631.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 627.7500 0.5200 627.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 623.7500 0.5200 623.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 619.7500 0.5200 619.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 615.7500 0.5200 615.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 611.7500 0.5200 611.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 607.7500 0.5200 607.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 603.7500 0.5200 603.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 599.7500 0.5200 599.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 595.7500 0.5200 595.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 591.7500 0.5200 591.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 587.7500 0.5200 587.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 583.7500 0.5200 583.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 579.7500 0.5200 579.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 575.7500 0.5200 575.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 571.7500 0.5200 571.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 567.7500 0.5200 567.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 563.7500 0.5200 563.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 559.7500 0.5200 559.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 555.7500 0.5200 555.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 551.7500 0.5200 551.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 547.7500 0.5200 547.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 543.7500 0.5200 543.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 539.7500 0.5200 539.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 535.7500 0.5200 535.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 531.7500 0.5200 531.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 527.7500 0.5200 527.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 523.7500 0.5200 523.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 519.7500 0.5200 519.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 515.7500 0.5200 515.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 511.7500 0.5200 511.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 507.7500 0.5200 507.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 503.7500 0.5200 503.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 499.7500 0.5200 499.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 495.7500 0.5200 495.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 491.7500 0.5200 491.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 487.7500 0.5200 487.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 483.7500 0.5200 483.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 479.7500 0.5200 479.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 475.7500 0.5200 475.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 471.7500 0.5200 471.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 444.1500 1420.0000 444.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 448.1500 1420.0000 448.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 452.1500 1420.0000 452.2500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 456.1500 1420.0000 456.2500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 460.1500 1420.0000 460.2500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 464.1500 1420.0000 464.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 468.1500 1420.0000 468.2500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 472.1500 1420.0000 472.2500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 476.1500 1420.0000 476.2500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 480.1500 1420.0000 480.2500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 484.1500 1420.0000 484.2500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 488.1500 1420.0000 488.2500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 492.1500 1420.0000 492.2500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 496.1500 1420.0000 496.2500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 500.1500 1420.0000 500.2500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 504.1500 1420.0000 504.2500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 508.1500 1420.0000 508.2500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 512.1500 1420.0000 512.2500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 516.1500 1420.0000 516.2500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 520.1500 1420.0000 520.2500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 524.1500 1420.0000 524.2500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 528.1500 1420.0000 528.2500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 532.1500 1420.0000 532.2500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 536.1500 1420.0000 536.2500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 540.1500 1420.0000 540.2500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 544.1500 1420.0000 544.2500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 548.1500 1420.0000 548.2500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 552.1500 1420.0000 552.2500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 556.1500 1420.0000 556.2500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 560.1500 1420.0000 560.2500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 564.1500 1420.0000 564.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 568.1500 1420.0000 568.2500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 572.1500 1420.0000 572.2500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 576.1500 1420.0000 576.2500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 580.1500 1420.0000 580.2500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 584.1500 1420.0000 584.2500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 588.1500 1420.0000 588.2500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 592.1500 1420.0000 592.2500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 596.1500 1420.0000 596.2500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 600.1500 1420.0000 600.2500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 604.1500 1420.0000 604.2500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 608.1500 1420.0000 608.2500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 612.1500 1420.0000 612.2500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 616.1500 1420.0000 616.2500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 620.1500 1420.0000 620.2500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 624.1500 1420.0000 624.2500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 628.1500 1420.0000 628.2500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 632.1500 1420.0000 632.2500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 636.1500 1420.0000 636.2500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 640.1500 1420.0000 640.2500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 644.1500 1420.0000 644.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 648.1500 1420.0000 648.2500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 652.1500 1420.0000 652.2500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 656.1500 1420.0000 656.2500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 660.1500 1420.0000 660.2500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 664.1500 1420.0000 664.2500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 668.1500 1420.0000 668.2500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 672.1500 1420.0000 672.2500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 676.1500 1420.0000 676.2500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 680.1500 1420.0000 680.2500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 684.1500 1420.0000 684.2500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 688.1500 1420.0000 688.2500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 692.1500 1420.0000 692.2500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 696.1500 1420.0000 696.2500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 700.1500 1420.0000 700.2500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 704.1500 1420.0000 704.2500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 708.1500 1420.0000 708.2500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 712.1500 1420.0000 712.2500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 716.1500 1420.0000 716.2500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 720.1500 1420.0000 720.2500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 724.1500 1420.0000 724.2500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 728.1500 1420.0000 728.2500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 732.1500 1420.0000 732.2500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 736.1500 1420.0000 736.2500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 740.1500 1420.0000 740.2500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 744.1500 1420.0000 744.2500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 748.1500 1420.0000 748.2500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 752.1500 1420.0000 752.2500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 756.1500 1420.0000 756.2500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 760.1500 1420.0000 760.2500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 860.1500 1420.0000 860.2500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 864.1500 1420.0000 864.2500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 868.1500 1420.0000 868.2500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 872.1500 1420.0000 872.2500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 876.1500 1420.0000 876.2500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 880.1500 1420.0000 880.2500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 884.1500 1420.0000 884.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 888.1500 1420.0000 888.2500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 892.1500 1420.0000 892.2500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 896.1500 1420.0000 896.2500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 900.1500 1420.0000 900.2500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 904.1500 1420.0000 904.2500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 908.1500 1420.0000 908.2500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 912.1500 1420.0000 912.2500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 916.1500 1420.0000 916.2500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 920.1500 1420.0000 920.2500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 924.1500 1420.0000 924.2500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 928.1500 1420.0000 928.2500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 932.1500 1420.0000 932.2500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 936.1500 1420.0000 936.2500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 940.1500 1420.0000 940.2500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 944.1500 1420.0000 944.2500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 948.1500 1420.0000 948.2500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 952.1500 1420.0000 952.2500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 956.1500 1420.0000 956.2500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 960.1500 1420.0000 960.2500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 964.1500 1420.0000 964.2500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 968.1500 1420.0000 968.2500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 972.1500 1420.0000 972.2500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 976.1500 1420.0000 976.2500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 980.1500 1420.0000 980.2500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 984.1500 1420.0000 984.2500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 988.1500 1420.0000 988.2500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 992.1500 1420.0000 992.2500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 996.1500 1420.0000 996.2500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1000.1500 1420.0000 1000.2500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1004.1500 1420.0000 1004.2500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1008.1500 1420.0000 1008.2500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1012.1500 1420.0000 1012.2500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1016.1500 1420.0000 1016.2500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1020.1500 1420.0000 1020.2500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1024.1500 1420.0000 1024.2500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1028.1500 1420.0000 1028.2500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1032.1500 1420.0000 1032.2500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1036.1500 1420.0000 1036.2500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1040.1500 1420.0000 1040.2500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1044.1500 1420.0000 1044.2500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1048.1500 1420.0000 1048.2500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1052.1500 1420.0000 1052.2500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1056.1500 1420.0000 1056.2500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1060.1500 1420.0000 1060.2500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1064.1500 1420.0000 1064.2500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1068.1500 1420.0000 1068.2500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1072.1500 1420.0000 1072.2500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1076.1500 1420.0000 1076.2500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1080.1500 1420.0000 1080.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1084.1500 1420.0000 1084.2500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1088.1500 1420.0000 1088.2500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1092.1500 1420.0000 1092.2500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1096.1500 1420.0000 1096.2500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1100.1500 1420.0000 1100.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1104.1500 1420.0000 1104.2500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1108.1500 1420.0000 1108.2500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1112.1500 1420.0000 1112.2500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1116.1500 1420.0000 1116.2500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1120.1500 1420.0000 1120.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1124.1500 1420.0000 1124.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1128.1500 1420.0000 1128.2500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1132.1500 1420.0000 1132.2500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1136.1500 1420.0000 1136.2500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1140.1500 1420.0000 1140.2500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1144.1500 1420.0000 1144.2500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1148.1500 1420.0000 1148.2500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1152.1500 1420.0000 1152.2500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1156.1500 1420.0000 1156.2500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1160.1500 1420.0000 1160.2500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1164.1500 1420.0000 1164.2500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1168.1500 1420.0000 1168.2500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1172.1500 1420.0000 1172.2500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1419.4800 1176.1500 1420.0000 1176.2500 ;
    END
  END out[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1015.7500 0.5200 1015.8500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1011.7500 0.5200 1011.8500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1007.7500 0.5200 1007.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1003.7500 0.5200 1003.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 999.7500 0.5200 999.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 995.7500 0.5200 995.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 991.7500 0.5200 991.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 987.7500 0.5200 987.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 983.7500 0.5200 983.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 459.7500 0.5200 459.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 455.7500 0.5200 455.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 451.7500 0.5200 451.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 447.7500 0.5200 447.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 443.7500 0.5200 443.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 439.7500 0.5200 439.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 435.7500 0.5200 435.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 431.7500 0.5200 431.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 427.7500 0.5200 427.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 423.7500 0.5200 423.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1059.7500 0.5200 1059.8500 ;
    END
  END reset
  PIN fifo_ext_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 467.7500 0.5200 467.8500 ;
    END
  END fifo_ext_rd
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
    LAYER M3 ;
      RECT 0.0000 809.9500 1420.0000 1620.0000 ;
      RECT 0.6200 809.6500 1420.0000 809.9500 ;
      RECT 0.0000 0.0000 1420.0000 809.6500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
    LAYER M5 ;
      RECT 0.0000 1176.3500 1420.0000 1620.0000 ;
      RECT 0.0000 1176.0500 1419.3800 1176.3500 ;
      RECT 0.0000 1172.3500 1420.0000 1176.0500 ;
      RECT 0.0000 1172.0500 1419.3800 1172.3500 ;
      RECT 0.0000 1168.3500 1420.0000 1172.0500 ;
      RECT 0.0000 1168.0500 1419.3800 1168.3500 ;
      RECT 0.0000 1164.3500 1420.0000 1168.0500 ;
      RECT 0.0000 1164.0500 1419.3800 1164.3500 ;
      RECT 0.0000 1160.3500 1420.0000 1164.0500 ;
      RECT 0.0000 1160.0500 1419.3800 1160.3500 ;
      RECT 0.0000 1156.3500 1420.0000 1160.0500 ;
      RECT 0.0000 1156.0500 1419.3800 1156.3500 ;
      RECT 0.0000 1155.9500 1420.0000 1156.0500 ;
      RECT 0.6200 1155.6500 1420.0000 1155.9500 ;
      RECT 0.0000 1152.3500 1420.0000 1155.6500 ;
      RECT 0.0000 1152.0500 1419.3800 1152.3500 ;
      RECT 0.0000 1151.9500 1420.0000 1152.0500 ;
      RECT 0.6200 1151.6500 1420.0000 1151.9500 ;
      RECT 0.0000 1148.3500 1420.0000 1151.6500 ;
      RECT 0.0000 1148.0500 1419.3800 1148.3500 ;
      RECT 0.0000 1147.9500 1420.0000 1148.0500 ;
      RECT 0.6200 1147.6500 1420.0000 1147.9500 ;
      RECT 0.0000 1144.3500 1420.0000 1147.6500 ;
      RECT 0.0000 1144.0500 1419.3800 1144.3500 ;
      RECT 0.0000 1143.9500 1420.0000 1144.0500 ;
      RECT 0.6200 1143.6500 1420.0000 1143.9500 ;
      RECT 0.0000 1140.3500 1420.0000 1143.6500 ;
      RECT 0.0000 1140.0500 1419.3800 1140.3500 ;
      RECT 0.0000 1139.9500 1420.0000 1140.0500 ;
      RECT 0.6200 1139.6500 1420.0000 1139.9500 ;
      RECT 0.0000 1136.3500 1420.0000 1139.6500 ;
      RECT 0.0000 1136.0500 1419.3800 1136.3500 ;
      RECT 0.0000 1135.9500 1420.0000 1136.0500 ;
      RECT 0.6200 1135.6500 1420.0000 1135.9500 ;
      RECT 0.0000 1132.3500 1420.0000 1135.6500 ;
      RECT 0.0000 1132.0500 1419.3800 1132.3500 ;
      RECT 0.0000 1131.9500 1420.0000 1132.0500 ;
      RECT 0.6200 1131.6500 1420.0000 1131.9500 ;
      RECT 0.0000 1128.3500 1420.0000 1131.6500 ;
      RECT 0.0000 1128.0500 1419.3800 1128.3500 ;
      RECT 0.0000 1127.9500 1420.0000 1128.0500 ;
      RECT 0.6200 1127.6500 1420.0000 1127.9500 ;
      RECT 0.0000 1124.3500 1420.0000 1127.6500 ;
      RECT 0.0000 1124.0500 1419.3800 1124.3500 ;
      RECT 0.0000 1123.9500 1420.0000 1124.0500 ;
      RECT 0.6200 1123.6500 1420.0000 1123.9500 ;
      RECT 0.0000 1120.3500 1420.0000 1123.6500 ;
      RECT 0.0000 1120.0500 1419.3800 1120.3500 ;
      RECT 0.0000 1119.9500 1420.0000 1120.0500 ;
      RECT 0.6200 1119.6500 1420.0000 1119.9500 ;
      RECT 0.0000 1116.3500 1420.0000 1119.6500 ;
      RECT 0.0000 1116.0500 1419.3800 1116.3500 ;
      RECT 0.0000 1115.9500 1420.0000 1116.0500 ;
      RECT 0.6200 1115.6500 1420.0000 1115.9500 ;
      RECT 0.0000 1112.3500 1420.0000 1115.6500 ;
      RECT 0.0000 1112.0500 1419.3800 1112.3500 ;
      RECT 0.0000 1111.9500 1420.0000 1112.0500 ;
      RECT 0.6200 1111.6500 1420.0000 1111.9500 ;
      RECT 0.0000 1108.3500 1420.0000 1111.6500 ;
      RECT 0.0000 1108.0500 1419.3800 1108.3500 ;
      RECT 0.0000 1107.9500 1420.0000 1108.0500 ;
      RECT 0.6200 1107.6500 1420.0000 1107.9500 ;
      RECT 0.0000 1104.3500 1420.0000 1107.6500 ;
      RECT 0.0000 1104.0500 1419.3800 1104.3500 ;
      RECT 0.0000 1103.9500 1420.0000 1104.0500 ;
      RECT 0.6200 1103.6500 1420.0000 1103.9500 ;
      RECT 0.0000 1100.3500 1420.0000 1103.6500 ;
      RECT 0.0000 1100.0500 1419.3800 1100.3500 ;
      RECT 0.0000 1099.9500 1420.0000 1100.0500 ;
      RECT 0.6200 1099.6500 1420.0000 1099.9500 ;
      RECT 0.0000 1096.3500 1420.0000 1099.6500 ;
      RECT 0.0000 1096.0500 1419.3800 1096.3500 ;
      RECT 0.0000 1095.9500 1420.0000 1096.0500 ;
      RECT 0.6200 1095.6500 1420.0000 1095.9500 ;
      RECT 0.0000 1092.3500 1420.0000 1095.6500 ;
      RECT 0.0000 1092.0500 1419.3800 1092.3500 ;
      RECT 0.0000 1091.9500 1420.0000 1092.0500 ;
      RECT 0.6200 1091.6500 1420.0000 1091.9500 ;
      RECT 0.0000 1088.3500 1420.0000 1091.6500 ;
      RECT 0.0000 1088.0500 1419.3800 1088.3500 ;
      RECT 0.0000 1087.9500 1420.0000 1088.0500 ;
      RECT 0.6200 1087.6500 1420.0000 1087.9500 ;
      RECT 0.0000 1084.3500 1420.0000 1087.6500 ;
      RECT 0.0000 1084.0500 1419.3800 1084.3500 ;
      RECT 0.0000 1083.9500 1420.0000 1084.0500 ;
      RECT 0.6200 1083.6500 1420.0000 1083.9500 ;
      RECT 0.0000 1080.3500 1420.0000 1083.6500 ;
      RECT 0.0000 1080.0500 1419.3800 1080.3500 ;
      RECT 0.0000 1079.9500 1420.0000 1080.0500 ;
      RECT 0.6200 1079.6500 1420.0000 1079.9500 ;
      RECT 0.0000 1076.3500 1420.0000 1079.6500 ;
      RECT 0.0000 1076.0500 1419.3800 1076.3500 ;
      RECT 0.0000 1075.9500 1420.0000 1076.0500 ;
      RECT 0.6200 1075.6500 1420.0000 1075.9500 ;
      RECT 0.0000 1072.3500 1420.0000 1075.6500 ;
      RECT 0.0000 1072.0500 1419.3800 1072.3500 ;
      RECT 0.0000 1071.9500 1420.0000 1072.0500 ;
      RECT 0.6200 1071.6500 1420.0000 1071.9500 ;
      RECT 0.0000 1068.3500 1420.0000 1071.6500 ;
      RECT 0.0000 1068.0500 1419.3800 1068.3500 ;
      RECT 0.0000 1067.9500 1420.0000 1068.0500 ;
      RECT 0.6200 1067.6500 1420.0000 1067.9500 ;
      RECT 0.0000 1064.3500 1420.0000 1067.6500 ;
      RECT 0.0000 1064.0500 1419.3800 1064.3500 ;
      RECT 0.0000 1063.9500 1420.0000 1064.0500 ;
      RECT 0.6200 1063.6500 1420.0000 1063.9500 ;
      RECT 0.0000 1060.3500 1420.0000 1063.6500 ;
      RECT 0.0000 1060.0500 1419.3800 1060.3500 ;
      RECT 0.0000 1059.9500 1420.0000 1060.0500 ;
      RECT 0.6200 1059.6500 1420.0000 1059.9500 ;
      RECT 0.0000 1056.3500 1420.0000 1059.6500 ;
      RECT 0.0000 1056.0500 1419.3800 1056.3500 ;
      RECT 0.0000 1052.3500 1420.0000 1056.0500 ;
      RECT 0.0000 1052.0500 1419.3800 1052.3500 ;
      RECT 0.0000 1048.3500 1420.0000 1052.0500 ;
      RECT 0.0000 1048.0500 1419.3800 1048.3500 ;
      RECT 0.0000 1044.3500 1420.0000 1048.0500 ;
      RECT 0.0000 1044.0500 1419.3800 1044.3500 ;
      RECT 0.0000 1040.3500 1420.0000 1044.0500 ;
      RECT 0.0000 1040.0500 1419.3800 1040.3500 ;
      RECT 0.0000 1036.3500 1420.0000 1040.0500 ;
      RECT 0.0000 1036.0500 1419.3800 1036.3500 ;
      RECT 0.0000 1032.3500 1420.0000 1036.0500 ;
      RECT 0.0000 1032.0500 1419.3800 1032.3500 ;
      RECT 0.0000 1028.3500 1420.0000 1032.0500 ;
      RECT 0.0000 1028.0500 1419.3800 1028.3500 ;
      RECT 0.0000 1024.3500 1420.0000 1028.0500 ;
      RECT 0.0000 1024.0500 1419.3800 1024.3500 ;
      RECT 0.0000 1020.3500 1420.0000 1024.0500 ;
      RECT 0.0000 1020.0500 1419.3800 1020.3500 ;
      RECT 0.0000 1016.3500 1420.0000 1020.0500 ;
      RECT 0.0000 1016.0500 1419.3800 1016.3500 ;
      RECT 0.0000 1015.9500 1420.0000 1016.0500 ;
      RECT 0.6200 1015.6500 1420.0000 1015.9500 ;
      RECT 0.0000 1012.3500 1420.0000 1015.6500 ;
      RECT 0.0000 1012.0500 1419.3800 1012.3500 ;
      RECT 0.0000 1011.9500 1420.0000 1012.0500 ;
      RECT 0.6200 1011.6500 1420.0000 1011.9500 ;
      RECT 0.0000 1008.3500 1420.0000 1011.6500 ;
      RECT 0.0000 1008.0500 1419.3800 1008.3500 ;
      RECT 0.0000 1007.9500 1420.0000 1008.0500 ;
      RECT 0.6200 1007.6500 1420.0000 1007.9500 ;
      RECT 0.0000 1004.3500 1420.0000 1007.6500 ;
      RECT 0.0000 1004.0500 1419.3800 1004.3500 ;
      RECT 0.0000 1003.9500 1420.0000 1004.0500 ;
      RECT 0.6200 1003.6500 1420.0000 1003.9500 ;
      RECT 0.0000 1000.3500 1420.0000 1003.6500 ;
      RECT 0.0000 1000.0500 1419.3800 1000.3500 ;
      RECT 0.0000 999.9500 1420.0000 1000.0500 ;
      RECT 0.6200 999.6500 1420.0000 999.9500 ;
      RECT 0.0000 996.3500 1420.0000 999.6500 ;
      RECT 0.0000 996.0500 1419.3800 996.3500 ;
      RECT 0.0000 995.9500 1420.0000 996.0500 ;
      RECT 0.6200 995.6500 1420.0000 995.9500 ;
      RECT 0.0000 992.3500 1420.0000 995.6500 ;
      RECT 0.0000 992.0500 1419.3800 992.3500 ;
      RECT 0.0000 991.9500 1420.0000 992.0500 ;
      RECT 0.6200 991.6500 1420.0000 991.9500 ;
      RECT 0.0000 988.3500 1420.0000 991.6500 ;
      RECT 0.0000 988.0500 1419.3800 988.3500 ;
      RECT 0.0000 987.9500 1420.0000 988.0500 ;
      RECT 0.6200 987.6500 1420.0000 987.9500 ;
      RECT 0.0000 984.3500 1420.0000 987.6500 ;
      RECT 0.0000 984.0500 1419.3800 984.3500 ;
      RECT 0.0000 983.9500 1420.0000 984.0500 ;
      RECT 0.6200 983.6500 1420.0000 983.9500 ;
      RECT 0.0000 980.3500 1420.0000 983.6500 ;
      RECT 0.0000 980.0500 1419.3800 980.3500 ;
      RECT 0.0000 979.9500 1420.0000 980.0500 ;
      RECT 0.6200 979.6500 1420.0000 979.9500 ;
      RECT 0.0000 976.3500 1420.0000 979.6500 ;
      RECT 0.0000 976.0500 1419.3800 976.3500 ;
      RECT 0.0000 975.9500 1420.0000 976.0500 ;
      RECT 0.6200 975.6500 1420.0000 975.9500 ;
      RECT 0.0000 972.3500 1420.0000 975.6500 ;
      RECT 0.0000 972.0500 1419.3800 972.3500 ;
      RECT 0.0000 971.9500 1420.0000 972.0500 ;
      RECT 0.6200 971.6500 1420.0000 971.9500 ;
      RECT 0.0000 968.3500 1420.0000 971.6500 ;
      RECT 0.0000 968.0500 1419.3800 968.3500 ;
      RECT 0.0000 967.9500 1420.0000 968.0500 ;
      RECT 0.6200 967.6500 1420.0000 967.9500 ;
      RECT 0.0000 964.3500 1420.0000 967.6500 ;
      RECT 0.0000 964.0500 1419.3800 964.3500 ;
      RECT 0.0000 963.9500 1420.0000 964.0500 ;
      RECT 0.6200 963.6500 1420.0000 963.9500 ;
      RECT 0.0000 960.3500 1420.0000 963.6500 ;
      RECT 0.0000 960.0500 1419.3800 960.3500 ;
      RECT 0.0000 959.9500 1420.0000 960.0500 ;
      RECT 0.6200 959.6500 1420.0000 959.9500 ;
      RECT 0.0000 956.3500 1420.0000 959.6500 ;
      RECT 0.0000 956.0500 1419.3800 956.3500 ;
      RECT 0.0000 955.9500 1420.0000 956.0500 ;
      RECT 0.6200 955.6500 1420.0000 955.9500 ;
      RECT 0.0000 952.3500 1420.0000 955.6500 ;
      RECT 0.0000 952.0500 1419.3800 952.3500 ;
      RECT 0.0000 951.9500 1420.0000 952.0500 ;
      RECT 0.6200 951.6500 1420.0000 951.9500 ;
      RECT 0.0000 948.3500 1420.0000 951.6500 ;
      RECT 0.0000 948.0500 1419.3800 948.3500 ;
      RECT 0.0000 947.9500 1420.0000 948.0500 ;
      RECT 0.6200 947.6500 1420.0000 947.9500 ;
      RECT 0.0000 944.3500 1420.0000 947.6500 ;
      RECT 0.0000 944.0500 1419.3800 944.3500 ;
      RECT 0.0000 943.9500 1420.0000 944.0500 ;
      RECT 0.6200 943.6500 1420.0000 943.9500 ;
      RECT 0.0000 940.3500 1420.0000 943.6500 ;
      RECT 0.0000 940.0500 1419.3800 940.3500 ;
      RECT 0.0000 939.9500 1420.0000 940.0500 ;
      RECT 0.6200 939.6500 1420.0000 939.9500 ;
      RECT 0.0000 936.3500 1420.0000 939.6500 ;
      RECT 0.0000 936.0500 1419.3800 936.3500 ;
      RECT 0.0000 935.9500 1420.0000 936.0500 ;
      RECT 0.6200 935.6500 1420.0000 935.9500 ;
      RECT 0.0000 932.3500 1420.0000 935.6500 ;
      RECT 0.0000 932.0500 1419.3800 932.3500 ;
      RECT 0.0000 931.9500 1420.0000 932.0500 ;
      RECT 0.6200 931.6500 1420.0000 931.9500 ;
      RECT 0.0000 928.3500 1420.0000 931.6500 ;
      RECT 0.0000 928.0500 1419.3800 928.3500 ;
      RECT 0.0000 927.9500 1420.0000 928.0500 ;
      RECT 0.6200 927.6500 1420.0000 927.9500 ;
      RECT 0.0000 924.3500 1420.0000 927.6500 ;
      RECT 0.0000 924.0500 1419.3800 924.3500 ;
      RECT 0.0000 923.9500 1420.0000 924.0500 ;
      RECT 0.6200 923.6500 1420.0000 923.9500 ;
      RECT 0.0000 920.3500 1420.0000 923.6500 ;
      RECT 0.0000 920.0500 1419.3800 920.3500 ;
      RECT 0.0000 919.9500 1420.0000 920.0500 ;
      RECT 0.6200 919.6500 1420.0000 919.9500 ;
      RECT 0.0000 916.3500 1420.0000 919.6500 ;
      RECT 0.0000 916.0500 1419.3800 916.3500 ;
      RECT 0.0000 915.9500 1420.0000 916.0500 ;
      RECT 0.6200 915.6500 1420.0000 915.9500 ;
      RECT 0.0000 912.3500 1420.0000 915.6500 ;
      RECT 0.0000 912.0500 1419.3800 912.3500 ;
      RECT 0.0000 911.9500 1420.0000 912.0500 ;
      RECT 0.6200 911.6500 1420.0000 911.9500 ;
      RECT 0.0000 908.3500 1420.0000 911.6500 ;
      RECT 0.0000 908.0500 1419.3800 908.3500 ;
      RECT 0.0000 907.9500 1420.0000 908.0500 ;
      RECT 0.6200 907.6500 1420.0000 907.9500 ;
      RECT 0.0000 904.3500 1420.0000 907.6500 ;
      RECT 0.0000 904.0500 1419.3800 904.3500 ;
      RECT 0.0000 903.9500 1420.0000 904.0500 ;
      RECT 0.6200 903.6500 1420.0000 903.9500 ;
      RECT 0.0000 900.3500 1420.0000 903.6500 ;
      RECT 0.0000 900.0500 1419.3800 900.3500 ;
      RECT 0.0000 899.9500 1420.0000 900.0500 ;
      RECT 0.6200 899.6500 1420.0000 899.9500 ;
      RECT 0.0000 896.3500 1420.0000 899.6500 ;
      RECT 0.0000 896.0500 1419.3800 896.3500 ;
      RECT 0.0000 895.9500 1420.0000 896.0500 ;
      RECT 0.6200 895.6500 1420.0000 895.9500 ;
      RECT 0.0000 892.3500 1420.0000 895.6500 ;
      RECT 0.0000 892.0500 1419.3800 892.3500 ;
      RECT 0.0000 891.9500 1420.0000 892.0500 ;
      RECT 0.6200 891.6500 1420.0000 891.9500 ;
      RECT 0.0000 888.3500 1420.0000 891.6500 ;
      RECT 0.0000 888.0500 1419.3800 888.3500 ;
      RECT 0.0000 887.9500 1420.0000 888.0500 ;
      RECT 0.6200 887.6500 1420.0000 887.9500 ;
      RECT 0.0000 884.3500 1420.0000 887.6500 ;
      RECT 0.0000 884.0500 1419.3800 884.3500 ;
      RECT 0.0000 883.9500 1420.0000 884.0500 ;
      RECT 0.6200 883.6500 1420.0000 883.9500 ;
      RECT 0.0000 880.3500 1420.0000 883.6500 ;
      RECT 0.0000 880.0500 1419.3800 880.3500 ;
      RECT 0.0000 879.9500 1420.0000 880.0500 ;
      RECT 0.6200 879.6500 1420.0000 879.9500 ;
      RECT 0.0000 876.3500 1420.0000 879.6500 ;
      RECT 0.0000 876.0500 1419.3800 876.3500 ;
      RECT 0.0000 875.9500 1420.0000 876.0500 ;
      RECT 0.6200 875.6500 1420.0000 875.9500 ;
      RECT 0.0000 872.3500 1420.0000 875.6500 ;
      RECT 0.0000 872.0500 1419.3800 872.3500 ;
      RECT 0.0000 871.9500 1420.0000 872.0500 ;
      RECT 0.6200 871.6500 1420.0000 871.9500 ;
      RECT 0.0000 868.3500 1420.0000 871.6500 ;
      RECT 0.0000 868.0500 1419.3800 868.3500 ;
      RECT 0.0000 867.9500 1420.0000 868.0500 ;
      RECT 0.6200 867.6500 1420.0000 867.9500 ;
      RECT 0.0000 864.3500 1420.0000 867.6500 ;
      RECT 0.0000 864.0500 1419.3800 864.3500 ;
      RECT 0.0000 863.9500 1420.0000 864.0500 ;
      RECT 0.6200 863.6500 1420.0000 863.9500 ;
      RECT 0.0000 860.3500 1420.0000 863.6500 ;
      RECT 0.0000 860.0500 1419.3800 860.3500 ;
      RECT 0.0000 859.9500 1420.0000 860.0500 ;
      RECT 0.6200 859.6500 1420.0000 859.9500 ;
      RECT 0.0000 856.3500 1420.0000 859.6500 ;
      RECT 0.0000 856.0500 1419.3800 856.3500 ;
      RECT 0.0000 855.9500 1420.0000 856.0500 ;
      RECT 0.6200 855.6500 1420.0000 855.9500 ;
      RECT 0.0000 852.3500 1420.0000 855.6500 ;
      RECT 0.0000 852.0500 1419.3800 852.3500 ;
      RECT 0.0000 851.9500 1420.0000 852.0500 ;
      RECT 0.6200 851.6500 1420.0000 851.9500 ;
      RECT 0.0000 848.3500 1420.0000 851.6500 ;
      RECT 0.0000 848.0500 1419.3800 848.3500 ;
      RECT 0.0000 847.9500 1420.0000 848.0500 ;
      RECT 0.6200 847.6500 1420.0000 847.9500 ;
      RECT 0.0000 844.3500 1420.0000 847.6500 ;
      RECT 0.0000 844.0500 1419.3800 844.3500 ;
      RECT 0.0000 843.9500 1420.0000 844.0500 ;
      RECT 0.6200 843.6500 1420.0000 843.9500 ;
      RECT 0.0000 840.3500 1420.0000 843.6500 ;
      RECT 0.0000 840.0500 1419.3800 840.3500 ;
      RECT 0.0000 839.9500 1420.0000 840.0500 ;
      RECT 0.6200 839.6500 1420.0000 839.9500 ;
      RECT 0.0000 836.3500 1420.0000 839.6500 ;
      RECT 0.0000 836.0500 1419.3800 836.3500 ;
      RECT 0.0000 835.9500 1420.0000 836.0500 ;
      RECT 0.6200 835.6500 1420.0000 835.9500 ;
      RECT 0.0000 832.3500 1420.0000 835.6500 ;
      RECT 0.0000 832.0500 1419.3800 832.3500 ;
      RECT 0.0000 831.9500 1420.0000 832.0500 ;
      RECT 0.6200 831.6500 1420.0000 831.9500 ;
      RECT 0.0000 828.3500 1420.0000 831.6500 ;
      RECT 0.0000 828.0500 1419.3800 828.3500 ;
      RECT 0.0000 827.9500 1420.0000 828.0500 ;
      RECT 0.6200 827.6500 1420.0000 827.9500 ;
      RECT 0.0000 824.3500 1420.0000 827.6500 ;
      RECT 0.0000 824.0500 1419.3800 824.3500 ;
      RECT 0.0000 823.9500 1420.0000 824.0500 ;
      RECT 0.6200 823.6500 1420.0000 823.9500 ;
      RECT 0.0000 820.3500 1420.0000 823.6500 ;
      RECT 0.0000 820.0500 1419.3800 820.3500 ;
      RECT 0.0000 819.9500 1420.0000 820.0500 ;
      RECT 0.6200 819.6500 1420.0000 819.9500 ;
      RECT 0.0000 816.3500 1420.0000 819.6500 ;
      RECT 0.0000 816.0500 1419.3800 816.3500 ;
      RECT 0.0000 815.9500 1420.0000 816.0500 ;
      RECT 0.6200 815.6500 1420.0000 815.9500 ;
      RECT 0.0000 812.3500 1420.0000 815.6500 ;
      RECT 0.0000 812.0500 1419.3800 812.3500 ;
      RECT 0.0000 811.9500 1420.0000 812.0500 ;
      RECT 0.6200 811.6500 1420.0000 811.9500 ;
      RECT 0.0000 808.3500 1420.0000 811.6500 ;
      RECT 0.0000 808.0500 1419.3800 808.3500 ;
      RECT 0.0000 807.9500 1420.0000 808.0500 ;
      RECT 0.6200 807.6500 1420.0000 807.9500 ;
      RECT 0.0000 804.3500 1420.0000 807.6500 ;
      RECT 0.0000 804.0500 1419.3800 804.3500 ;
      RECT 0.0000 803.9500 1420.0000 804.0500 ;
      RECT 0.6200 803.6500 1420.0000 803.9500 ;
      RECT 0.0000 800.3500 1420.0000 803.6500 ;
      RECT 0.0000 800.0500 1419.3800 800.3500 ;
      RECT 0.0000 799.9500 1420.0000 800.0500 ;
      RECT 0.6200 799.6500 1420.0000 799.9500 ;
      RECT 0.0000 796.3500 1420.0000 799.6500 ;
      RECT 0.0000 796.0500 1419.3800 796.3500 ;
      RECT 0.0000 795.9500 1420.0000 796.0500 ;
      RECT 0.6200 795.6500 1420.0000 795.9500 ;
      RECT 0.0000 792.3500 1420.0000 795.6500 ;
      RECT 0.0000 792.0500 1419.3800 792.3500 ;
      RECT 0.0000 791.9500 1420.0000 792.0500 ;
      RECT 0.6200 791.6500 1420.0000 791.9500 ;
      RECT 0.0000 788.3500 1420.0000 791.6500 ;
      RECT 0.0000 788.0500 1419.3800 788.3500 ;
      RECT 0.0000 787.9500 1420.0000 788.0500 ;
      RECT 0.6200 787.6500 1420.0000 787.9500 ;
      RECT 0.0000 784.3500 1420.0000 787.6500 ;
      RECT 0.0000 784.0500 1419.3800 784.3500 ;
      RECT 0.0000 783.9500 1420.0000 784.0500 ;
      RECT 0.6200 783.6500 1420.0000 783.9500 ;
      RECT 0.0000 780.3500 1420.0000 783.6500 ;
      RECT 0.0000 780.0500 1419.3800 780.3500 ;
      RECT 0.0000 779.9500 1420.0000 780.0500 ;
      RECT 0.6200 779.6500 1420.0000 779.9500 ;
      RECT 0.0000 776.3500 1420.0000 779.6500 ;
      RECT 0.0000 776.0500 1419.3800 776.3500 ;
      RECT 0.0000 775.9500 1420.0000 776.0500 ;
      RECT 0.6200 775.6500 1420.0000 775.9500 ;
      RECT 0.0000 772.3500 1420.0000 775.6500 ;
      RECT 0.0000 772.0500 1419.3800 772.3500 ;
      RECT 0.0000 771.9500 1420.0000 772.0500 ;
      RECT 0.6200 771.6500 1420.0000 771.9500 ;
      RECT 0.0000 768.3500 1420.0000 771.6500 ;
      RECT 0.0000 768.0500 1419.3800 768.3500 ;
      RECT 0.0000 767.9500 1420.0000 768.0500 ;
      RECT 0.6200 767.6500 1420.0000 767.9500 ;
      RECT 0.0000 764.3500 1420.0000 767.6500 ;
      RECT 0.0000 764.0500 1419.3800 764.3500 ;
      RECT 0.0000 763.9500 1420.0000 764.0500 ;
      RECT 0.6200 763.6500 1420.0000 763.9500 ;
      RECT 0.0000 760.3500 1420.0000 763.6500 ;
      RECT 0.0000 760.0500 1419.3800 760.3500 ;
      RECT 0.0000 759.9500 1420.0000 760.0500 ;
      RECT 0.6200 759.6500 1420.0000 759.9500 ;
      RECT 0.0000 756.3500 1420.0000 759.6500 ;
      RECT 0.0000 756.0500 1419.3800 756.3500 ;
      RECT 0.0000 755.9500 1420.0000 756.0500 ;
      RECT 0.6200 755.6500 1420.0000 755.9500 ;
      RECT 0.0000 752.3500 1420.0000 755.6500 ;
      RECT 0.0000 752.0500 1419.3800 752.3500 ;
      RECT 0.0000 751.9500 1420.0000 752.0500 ;
      RECT 0.6200 751.6500 1420.0000 751.9500 ;
      RECT 0.0000 748.3500 1420.0000 751.6500 ;
      RECT 0.0000 748.0500 1419.3800 748.3500 ;
      RECT 0.0000 747.9500 1420.0000 748.0500 ;
      RECT 0.6200 747.6500 1420.0000 747.9500 ;
      RECT 0.0000 744.3500 1420.0000 747.6500 ;
      RECT 0.0000 744.0500 1419.3800 744.3500 ;
      RECT 0.0000 743.9500 1420.0000 744.0500 ;
      RECT 0.6200 743.6500 1420.0000 743.9500 ;
      RECT 0.0000 740.3500 1420.0000 743.6500 ;
      RECT 0.0000 740.0500 1419.3800 740.3500 ;
      RECT 0.0000 739.9500 1420.0000 740.0500 ;
      RECT 0.6200 739.6500 1420.0000 739.9500 ;
      RECT 0.0000 736.3500 1420.0000 739.6500 ;
      RECT 0.0000 736.0500 1419.3800 736.3500 ;
      RECT 0.0000 735.9500 1420.0000 736.0500 ;
      RECT 0.6200 735.6500 1420.0000 735.9500 ;
      RECT 0.0000 732.3500 1420.0000 735.6500 ;
      RECT 0.0000 732.0500 1419.3800 732.3500 ;
      RECT 0.0000 731.9500 1420.0000 732.0500 ;
      RECT 0.6200 731.6500 1420.0000 731.9500 ;
      RECT 0.0000 728.3500 1420.0000 731.6500 ;
      RECT 0.0000 728.0500 1419.3800 728.3500 ;
      RECT 0.0000 727.9500 1420.0000 728.0500 ;
      RECT 0.6200 727.6500 1420.0000 727.9500 ;
      RECT 0.0000 724.3500 1420.0000 727.6500 ;
      RECT 0.0000 724.0500 1419.3800 724.3500 ;
      RECT 0.0000 723.9500 1420.0000 724.0500 ;
      RECT 0.6200 723.6500 1420.0000 723.9500 ;
      RECT 0.0000 720.3500 1420.0000 723.6500 ;
      RECT 0.0000 720.0500 1419.3800 720.3500 ;
      RECT 0.0000 719.9500 1420.0000 720.0500 ;
      RECT 0.6200 719.6500 1420.0000 719.9500 ;
      RECT 0.0000 716.3500 1420.0000 719.6500 ;
      RECT 0.0000 716.0500 1419.3800 716.3500 ;
      RECT 0.0000 715.9500 1420.0000 716.0500 ;
      RECT 0.6200 715.6500 1420.0000 715.9500 ;
      RECT 0.0000 712.3500 1420.0000 715.6500 ;
      RECT 0.0000 712.0500 1419.3800 712.3500 ;
      RECT 0.0000 711.9500 1420.0000 712.0500 ;
      RECT 0.6200 711.6500 1420.0000 711.9500 ;
      RECT 0.0000 708.3500 1420.0000 711.6500 ;
      RECT 0.0000 708.0500 1419.3800 708.3500 ;
      RECT 0.0000 707.9500 1420.0000 708.0500 ;
      RECT 0.6200 707.6500 1420.0000 707.9500 ;
      RECT 0.0000 704.3500 1420.0000 707.6500 ;
      RECT 0.0000 704.0500 1419.3800 704.3500 ;
      RECT 0.0000 703.9500 1420.0000 704.0500 ;
      RECT 0.6200 703.6500 1420.0000 703.9500 ;
      RECT 0.0000 700.3500 1420.0000 703.6500 ;
      RECT 0.0000 700.0500 1419.3800 700.3500 ;
      RECT 0.0000 699.9500 1420.0000 700.0500 ;
      RECT 0.6200 699.6500 1420.0000 699.9500 ;
      RECT 0.0000 696.3500 1420.0000 699.6500 ;
      RECT 0.0000 696.0500 1419.3800 696.3500 ;
      RECT 0.0000 695.9500 1420.0000 696.0500 ;
      RECT 0.6200 695.6500 1420.0000 695.9500 ;
      RECT 0.0000 692.3500 1420.0000 695.6500 ;
      RECT 0.0000 692.0500 1419.3800 692.3500 ;
      RECT 0.0000 691.9500 1420.0000 692.0500 ;
      RECT 0.6200 691.6500 1420.0000 691.9500 ;
      RECT 0.0000 688.3500 1420.0000 691.6500 ;
      RECT 0.0000 688.0500 1419.3800 688.3500 ;
      RECT 0.0000 687.9500 1420.0000 688.0500 ;
      RECT 0.6200 687.6500 1420.0000 687.9500 ;
      RECT 0.0000 684.3500 1420.0000 687.6500 ;
      RECT 0.0000 684.0500 1419.3800 684.3500 ;
      RECT 0.0000 683.9500 1420.0000 684.0500 ;
      RECT 0.6200 683.6500 1420.0000 683.9500 ;
      RECT 0.0000 680.3500 1420.0000 683.6500 ;
      RECT 0.0000 680.0500 1419.3800 680.3500 ;
      RECT 0.0000 679.9500 1420.0000 680.0500 ;
      RECT 0.6200 679.6500 1420.0000 679.9500 ;
      RECT 0.0000 676.3500 1420.0000 679.6500 ;
      RECT 0.0000 676.0500 1419.3800 676.3500 ;
      RECT 0.0000 675.9500 1420.0000 676.0500 ;
      RECT 0.6200 675.6500 1420.0000 675.9500 ;
      RECT 0.0000 672.3500 1420.0000 675.6500 ;
      RECT 0.0000 672.0500 1419.3800 672.3500 ;
      RECT 0.0000 671.9500 1420.0000 672.0500 ;
      RECT 0.6200 671.6500 1420.0000 671.9500 ;
      RECT 0.0000 668.3500 1420.0000 671.6500 ;
      RECT 0.0000 668.0500 1419.3800 668.3500 ;
      RECT 0.0000 667.9500 1420.0000 668.0500 ;
      RECT 0.6200 667.6500 1420.0000 667.9500 ;
      RECT 0.0000 664.3500 1420.0000 667.6500 ;
      RECT 0.0000 664.0500 1419.3800 664.3500 ;
      RECT 0.0000 663.9500 1420.0000 664.0500 ;
      RECT 0.6200 663.6500 1420.0000 663.9500 ;
      RECT 0.0000 660.3500 1420.0000 663.6500 ;
      RECT 0.0000 660.0500 1419.3800 660.3500 ;
      RECT 0.0000 659.9500 1420.0000 660.0500 ;
      RECT 0.6200 659.6500 1420.0000 659.9500 ;
      RECT 0.0000 656.3500 1420.0000 659.6500 ;
      RECT 0.0000 656.0500 1419.3800 656.3500 ;
      RECT 0.0000 655.9500 1420.0000 656.0500 ;
      RECT 0.6200 655.6500 1420.0000 655.9500 ;
      RECT 0.0000 652.3500 1420.0000 655.6500 ;
      RECT 0.0000 652.0500 1419.3800 652.3500 ;
      RECT 0.0000 651.9500 1420.0000 652.0500 ;
      RECT 0.6200 651.6500 1420.0000 651.9500 ;
      RECT 0.0000 648.3500 1420.0000 651.6500 ;
      RECT 0.0000 648.0500 1419.3800 648.3500 ;
      RECT 0.0000 647.9500 1420.0000 648.0500 ;
      RECT 0.6200 647.6500 1420.0000 647.9500 ;
      RECT 0.0000 644.3500 1420.0000 647.6500 ;
      RECT 0.0000 644.0500 1419.3800 644.3500 ;
      RECT 0.0000 643.9500 1420.0000 644.0500 ;
      RECT 0.6200 643.6500 1420.0000 643.9500 ;
      RECT 0.0000 640.3500 1420.0000 643.6500 ;
      RECT 0.0000 640.0500 1419.3800 640.3500 ;
      RECT 0.0000 639.9500 1420.0000 640.0500 ;
      RECT 0.6200 639.6500 1420.0000 639.9500 ;
      RECT 0.0000 636.3500 1420.0000 639.6500 ;
      RECT 0.0000 636.0500 1419.3800 636.3500 ;
      RECT 0.0000 635.9500 1420.0000 636.0500 ;
      RECT 0.6200 635.6500 1420.0000 635.9500 ;
      RECT 0.0000 632.3500 1420.0000 635.6500 ;
      RECT 0.0000 632.0500 1419.3800 632.3500 ;
      RECT 0.0000 631.9500 1420.0000 632.0500 ;
      RECT 0.6200 631.6500 1420.0000 631.9500 ;
      RECT 0.0000 628.3500 1420.0000 631.6500 ;
      RECT 0.0000 628.0500 1419.3800 628.3500 ;
      RECT 0.0000 627.9500 1420.0000 628.0500 ;
      RECT 0.6200 627.6500 1420.0000 627.9500 ;
      RECT 0.0000 624.3500 1420.0000 627.6500 ;
      RECT 0.0000 624.0500 1419.3800 624.3500 ;
      RECT 0.0000 623.9500 1420.0000 624.0500 ;
      RECT 0.6200 623.6500 1420.0000 623.9500 ;
      RECT 0.0000 620.3500 1420.0000 623.6500 ;
      RECT 0.0000 620.0500 1419.3800 620.3500 ;
      RECT 0.0000 619.9500 1420.0000 620.0500 ;
      RECT 0.6200 619.6500 1420.0000 619.9500 ;
      RECT 0.0000 616.3500 1420.0000 619.6500 ;
      RECT 0.0000 616.0500 1419.3800 616.3500 ;
      RECT 0.0000 615.9500 1420.0000 616.0500 ;
      RECT 0.6200 615.6500 1420.0000 615.9500 ;
      RECT 0.0000 612.3500 1420.0000 615.6500 ;
      RECT 0.0000 612.0500 1419.3800 612.3500 ;
      RECT 0.0000 611.9500 1420.0000 612.0500 ;
      RECT 0.6200 611.6500 1420.0000 611.9500 ;
      RECT 0.0000 608.3500 1420.0000 611.6500 ;
      RECT 0.0000 608.0500 1419.3800 608.3500 ;
      RECT 0.0000 607.9500 1420.0000 608.0500 ;
      RECT 0.6200 607.6500 1420.0000 607.9500 ;
      RECT 0.0000 604.3500 1420.0000 607.6500 ;
      RECT 0.0000 604.0500 1419.3800 604.3500 ;
      RECT 0.0000 603.9500 1420.0000 604.0500 ;
      RECT 0.6200 603.6500 1420.0000 603.9500 ;
      RECT 0.0000 600.3500 1420.0000 603.6500 ;
      RECT 0.0000 600.0500 1419.3800 600.3500 ;
      RECT 0.0000 599.9500 1420.0000 600.0500 ;
      RECT 0.6200 599.6500 1420.0000 599.9500 ;
      RECT 0.0000 596.3500 1420.0000 599.6500 ;
      RECT 0.0000 596.0500 1419.3800 596.3500 ;
      RECT 0.0000 595.9500 1420.0000 596.0500 ;
      RECT 0.6200 595.6500 1420.0000 595.9500 ;
      RECT 0.0000 592.3500 1420.0000 595.6500 ;
      RECT 0.0000 592.0500 1419.3800 592.3500 ;
      RECT 0.0000 591.9500 1420.0000 592.0500 ;
      RECT 0.6200 591.6500 1420.0000 591.9500 ;
      RECT 0.0000 588.3500 1420.0000 591.6500 ;
      RECT 0.0000 588.0500 1419.3800 588.3500 ;
      RECT 0.0000 587.9500 1420.0000 588.0500 ;
      RECT 0.6200 587.6500 1420.0000 587.9500 ;
      RECT 0.0000 584.3500 1420.0000 587.6500 ;
      RECT 0.0000 584.0500 1419.3800 584.3500 ;
      RECT 0.0000 583.9500 1420.0000 584.0500 ;
      RECT 0.6200 583.6500 1420.0000 583.9500 ;
      RECT 0.0000 580.3500 1420.0000 583.6500 ;
      RECT 0.0000 580.0500 1419.3800 580.3500 ;
      RECT 0.0000 579.9500 1420.0000 580.0500 ;
      RECT 0.6200 579.6500 1420.0000 579.9500 ;
      RECT 0.0000 576.3500 1420.0000 579.6500 ;
      RECT 0.0000 576.0500 1419.3800 576.3500 ;
      RECT 0.0000 575.9500 1420.0000 576.0500 ;
      RECT 0.6200 575.6500 1420.0000 575.9500 ;
      RECT 0.0000 572.3500 1420.0000 575.6500 ;
      RECT 0.0000 572.0500 1419.3800 572.3500 ;
      RECT 0.0000 571.9500 1420.0000 572.0500 ;
      RECT 0.6200 571.6500 1420.0000 571.9500 ;
      RECT 0.0000 568.3500 1420.0000 571.6500 ;
      RECT 0.0000 568.0500 1419.3800 568.3500 ;
      RECT 0.0000 567.9500 1420.0000 568.0500 ;
      RECT 0.6200 567.6500 1420.0000 567.9500 ;
      RECT 0.0000 564.3500 1420.0000 567.6500 ;
      RECT 0.0000 564.0500 1419.3800 564.3500 ;
      RECT 0.0000 563.9500 1420.0000 564.0500 ;
      RECT 0.6200 563.6500 1420.0000 563.9500 ;
      RECT 0.0000 560.3500 1420.0000 563.6500 ;
      RECT 0.0000 560.0500 1419.3800 560.3500 ;
      RECT 0.0000 559.9500 1420.0000 560.0500 ;
      RECT 0.6200 559.6500 1420.0000 559.9500 ;
      RECT 0.0000 556.3500 1420.0000 559.6500 ;
      RECT 0.0000 556.0500 1419.3800 556.3500 ;
      RECT 0.0000 555.9500 1420.0000 556.0500 ;
      RECT 0.6200 555.6500 1420.0000 555.9500 ;
      RECT 0.0000 552.3500 1420.0000 555.6500 ;
      RECT 0.0000 552.0500 1419.3800 552.3500 ;
      RECT 0.0000 551.9500 1420.0000 552.0500 ;
      RECT 0.6200 551.6500 1420.0000 551.9500 ;
      RECT 0.0000 548.3500 1420.0000 551.6500 ;
      RECT 0.0000 548.0500 1419.3800 548.3500 ;
      RECT 0.0000 547.9500 1420.0000 548.0500 ;
      RECT 0.6200 547.6500 1420.0000 547.9500 ;
      RECT 0.0000 544.3500 1420.0000 547.6500 ;
      RECT 0.0000 544.0500 1419.3800 544.3500 ;
      RECT 0.0000 543.9500 1420.0000 544.0500 ;
      RECT 0.6200 543.6500 1420.0000 543.9500 ;
      RECT 0.0000 540.3500 1420.0000 543.6500 ;
      RECT 0.0000 540.0500 1419.3800 540.3500 ;
      RECT 0.0000 539.9500 1420.0000 540.0500 ;
      RECT 0.6200 539.6500 1420.0000 539.9500 ;
      RECT 0.0000 536.3500 1420.0000 539.6500 ;
      RECT 0.0000 536.0500 1419.3800 536.3500 ;
      RECT 0.0000 535.9500 1420.0000 536.0500 ;
      RECT 0.6200 535.6500 1420.0000 535.9500 ;
      RECT 0.0000 532.3500 1420.0000 535.6500 ;
      RECT 0.0000 532.0500 1419.3800 532.3500 ;
      RECT 0.0000 531.9500 1420.0000 532.0500 ;
      RECT 0.6200 531.6500 1420.0000 531.9500 ;
      RECT 0.0000 528.3500 1420.0000 531.6500 ;
      RECT 0.0000 528.0500 1419.3800 528.3500 ;
      RECT 0.0000 527.9500 1420.0000 528.0500 ;
      RECT 0.6200 527.6500 1420.0000 527.9500 ;
      RECT 0.0000 524.3500 1420.0000 527.6500 ;
      RECT 0.0000 524.0500 1419.3800 524.3500 ;
      RECT 0.0000 523.9500 1420.0000 524.0500 ;
      RECT 0.6200 523.6500 1420.0000 523.9500 ;
      RECT 0.0000 520.3500 1420.0000 523.6500 ;
      RECT 0.0000 520.0500 1419.3800 520.3500 ;
      RECT 0.0000 519.9500 1420.0000 520.0500 ;
      RECT 0.6200 519.6500 1420.0000 519.9500 ;
      RECT 0.0000 516.3500 1420.0000 519.6500 ;
      RECT 0.0000 516.0500 1419.3800 516.3500 ;
      RECT 0.0000 515.9500 1420.0000 516.0500 ;
      RECT 0.6200 515.6500 1420.0000 515.9500 ;
      RECT 0.0000 512.3500 1420.0000 515.6500 ;
      RECT 0.0000 512.0500 1419.3800 512.3500 ;
      RECT 0.0000 511.9500 1420.0000 512.0500 ;
      RECT 0.6200 511.6500 1420.0000 511.9500 ;
      RECT 0.0000 508.3500 1420.0000 511.6500 ;
      RECT 0.0000 508.0500 1419.3800 508.3500 ;
      RECT 0.0000 507.9500 1420.0000 508.0500 ;
      RECT 0.6200 507.6500 1420.0000 507.9500 ;
      RECT 0.0000 504.3500 1420.0000 507.6500 ;
      RECT 0.0000 504.0500 1419.3800 504.3500 ;
      RECT 0.0000 503.9500 1420.0000 504.0500 ;
      RECT 0.6200 503.6500 1420.0000 503.9500 ;
      RECT 0.0000 500.3500 1420.0000 503.6500 ;
      RECT 0.0000 500.0500 1419.3800 500.3500 ;
      RECT 0.0000 499.9500 1420.0000 500.0500 ;
      RECT 0.6200 499.6500 1420.0000 499.9500 ;
      RECT 0.0000 496.3500 1420.0000 499.6500 ;
      RECT 0.0000 496.0500 1419.3800 496.3500 ;
      RECT 0.0000 495.9500 1420.0000 496.0500 ;
      RECT 0.6200 495.6500 1420.0000 495.9500 ;
      RECT 0.0000 492.3500 1420.0000 495.6500 ;
      RECT 0.0000 492.0500 1419.3800 492.3500 ;
      RECT 0.0000 491.9500 1420.0000 492.0500 ;
      RECT 0.6200 491.6500 1420.0000 491.9500 ;
      RECT 0.0000 488.3500 1420.0000 491.6500 ;
      RECT 0.0000 488.0500 1419.3800 488.3500 ;
      RECT 0.0000 487.9500 1420.0000 488.0500 ;
      RECT 0.6200 487.6500 1420.0000 487.9500 ;
      RECT 0.0000 484.3500 1420.0000 487.6500 ;
      RECT 0.0000 484.0500 1419.3800 484.3500 ;
      RECT 0.0000 483.9500 1420.0000 484.0500 ;
      RECT 0.6200 483.6500 1420.0000 483.9500 ;
      RECT 0.0000 480.3500 1420.0000 483.6500 ;
      RECT 0.0000 480.0500 1419.3800 480.3500 ;
      RECT 0.0000 479.9500 1420.0000 480.0500 ;
      RECT 0.6200 479.6500 1420.0000 479.9500 ;
      RECT 0.0000 476.3500 1420.0000 479.6500 ;
      RECT 0.0000 476.0500 1419.3800 476.3500 ;
      RECT 0.0000 475.9500 1420.0000 476.0500 ;
      RECT 0.6200 475.6500 1420.0000 475.9500 ;
      RECT 0.0000 472.3500 1420.0000 475.6500 ;
      RECT 0.0000 472.0500 1419.3800 472.3500 ;
      RECT 0.0000 471.9500 1420.0000 472.0500 ;
      RECT 0.6200 471.6500 1420.0000 471.9500 ;
      RECT 0.0000 468.3500 1420.0000 471.6500 ;
      RECT 0.0000 468.0500 1419.3800 468.3500 ;
      RECT 0.0000 467.9500 1420.0000 468.0500 ;
      RECT 0.6200 467.6500 1420.0000 467.9500 ;
      RECT 0.0000 464.3500 1420.0000 467.6500 ;
      RECT 0.0000 464.0500 1419.3800 464.3500 ;
      RECT 0.0000 460.3500 1420.0000 464.0500 ;
      RECT 0.0000 460.0500 1419.3800 460.3500 ;
      RECT 0.0000 459.9500 1420.0000 460.0500 ;
      RECT 0.6200 459.6500 1420.0000 459.9500 ;
      RECT 0.0000 456.3500 1420.0000 459.6500 ;
      RECT 0.0000 456.0500 1419.3800 456.3500 ;
      RECT 0.0000 455.9500 1420.0000 456.0500 ;
      RECT 0.6200 455.6500 1420.0000 455.9500 ;
      RECT 0.0000 452.3500 1420.0000 455.6500 ;
      RECT 0.0000 452.0500 1419.3800 452.3500 ;
      RECT 0.0000 451.9500 1420.0000 452.0500 ;
      RECT 0.6200 451.6500 1420.0000 451.9500 ;
      RECT 0.0000 448.3500 1420.0000 451.6500 ;
      RECT 0.0000 448.0500 1419.3800 448.3500 ;
      RECT 0.0000 447.9500 1420.0000 448.0500 ;
      RECT 0.6200 447.6500 1420.0000 447.9500 ;
      RECT 0.0000 444.3500 1420.0000 447.6500 ;
      RECT 0.0000 444.0500 1419.3800 444.3500 ;
      RECT 0.0000 443.9500 1420.0000 444.0500 ;
      RECT 0.6200 443.6500 1420.0000 443.9500 ;
      RECT 0.0000 439.9500 1420.0000 443.6500 ;
      RECT 0.6200 439.6500 1420.0000 439.9500 ;
      RECT 0.0000 435.9500 1420.0000 439.6500 ;
      RECT 0.6200 435.6500 1420.0000 435.9500 ;
      RECT 0.0000 431.9500 1420.0000 435.6500 ;
      RECT 0.6200 431.6500 1420.0000 431.9500 ;
      RECT 0.0000 427.9500 1420.0000 431.6500 ;
      RECT 0.6200 427.6500 1420.0000 427.9500 ;
      RECT 0.0000 423.9500 1420.0000 427.6500 ;
      RECT 0.6200 423.6500 1420.0000 423.9500 ;
      RECT 0.0000 0.0000 1420.0000 423.6500 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1420.0000 1620.0000 ;
  END
END core

END LIBRARY
