/home/linux/ieng6/ee260bwi25/jmsin/ece260_project/step3/pnr_fullchip/subckt/sram_w16.lef