##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Wed Mar 19 13:34:46 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1020.0000 BY 1620.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 463.7500 0.5200 463.8500 ;
    END
  END clk
  PIN sum_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1155.7500 0.5200 1155.8500 ;
    END
  END sum_in[23]
  PIN sum_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1151.7500 0.5200 1151.8500 ;
    END
  END sum_in[22]
  PIN sum_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1147.7500 0.5200 1147.8500 ;
    END
  END sum_in[21]
  PIN sum_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1143.7500 0.5200 1143.8500 ;
    END
  END sum_in[20]
  PIN sum_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1139.7500 0.5200 1139.8500 ;
    END
  END sum_in[19]
  PIN sum_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1135.7500 0.5200 1135.8500 ;
    END
  END sum_in[18]
  PIN sum_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1131.7500 0.5200 1131.8500 ;
    END
  END sum_in[17]
  PIN sum_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1127.7500 0.5200 1127.8500 ;
    END
  END sum_in[16]
  PIN sum_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1123.7500 0.5200 1123.8500 ;
    END
  END sum_in[15]
  PIN sum_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1119.7500 0.5200 1119.8500 ;
    END
  END sum_in[14]
  PIN sum_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1115.7500 0.5200 1115.8500 ;
    END
  END sum_in[13]
  PIN sum_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1111.7500 0.5200 1111.8500 ;
    END
  END sum_in[12]
  PIN sum_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1107.7500 0.5200 1107.8500 ;
    END
  END sum_in[11]
  PIN sum_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1103.7500 0.5200 1103.8500 ;
    END
  END sum_in[10]
  PIN sum_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1099.7500 0.5200 1099.8500 ;
    END
  END sum_in[9]
  PIN sum_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1095.7500 0.5200 1095.8500 ;
    END
  END sum_in[8]
  PIN sum_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1091.7500 0.5200 1091.8500 ;
    END
  END sum_in[7]
  PIN sum_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1087.7500 0.5200 1087.8500 ;
    END
  END sum_in[6]
  PIN sum_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1083.7500 0.5200 1083.8500 ;
    END
  END sum_in[5]
  PIN sum_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1079.7500 0.5200 1079.8500 ;
    END
  END sum_in[4]
  PIN sum_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1075.7500 0.5200 1075.8500 ;
    END
  END sum_in[3]
  PIN sum_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1071.7500 0.5200 1071.8500 ;
    END
  END sum_in[2]
  PIN sum_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1067.7500 0.5200 1067.8500 ;
    END
  END sum_in[1]
  PIN sum_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1063.7500 0.5200 1063.8500 ;
    END
  END sum_in[0]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1084.1500 1020.0000 1084.2500 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1088.1500 1020.0000 1088.2500 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1092.1500 1020.0000 1092.2500 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1096.1500 1020.0000 1096.2500 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1100.1500 1020.0000 1100.2500 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1104.1500 1020.0000 1104.2500 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1108.1500 1020.0000 1108.2500 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1112.1500 1020.0000 1112.2500 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1116.1500 1020.0000 1116.2500 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1120.1500 1020.0000 1120.2500 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1124.1500 1020.0000 1124.2500 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1128.1500 1020.0000 1128.2500 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1132.1500 1020.0000 1132.2500 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1136.1500 1020.0000 1136.2500 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1140.1500 1020.0000 1140.2500 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1144.1500 1020.0000 1144.2500 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1148.1500 1020.0000 1148.2500 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1152.1500 1020.0000 1152.2500 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1156.1500 1020.0000 1156.2500 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1160.1500 1020.0000 1160.2500 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1164.1500 1020.0000 1164.2500 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1168.1500 1020.0000 1168.2500 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1172.1500 1020.0000 1172.2500 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1176.1500 1020.0000 1176.2500 ;
    END
  END sum_out[0]
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1055.7500 0.5200 1055.8500 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1051.7500 0.5200 1051.8500 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1047.7500 0.5200 1047.8500 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1043.7500 0.5200 1043.8500 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1039.7500 0.5200 1039.8500 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1035.7500 0.5200 1035.8500 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1031.7500 0.5200 1031.8500 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1027.7500 0.5200 1027.8500 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1023.7500 0.5200 1023.8500 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1019.7500 0.5200 1019.8500 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1015.7500 0.5200 1015.8500 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1011.7500 0.5200 1011.8500 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1007.7500 0.5200 1007.8500 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1003.7500 0.5200 1003.8500 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 999.7500 0.5200 999.8500 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 995.7500 0.5200 995.8500 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 991.7500 0.5200 991.8500 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 987.7500 0.5200 987.8500 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 983.7500 0.5200 983.8500 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 979.7500 0.5200 979.8500 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 975.7500 0.5200 975.8500 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 971.7500 0.5200 971.8500 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 967.7500 0.5200 967.8500 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 963.7500 0.5200 963.8500 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 959.7500 0.5200 959.8500 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 955.7500 0.5200 955.8500 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 951.7500 0.5200 951.8500 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 947.7500 0.5200 947.8500 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 943.7500 0.5200 943.8500 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 939.7500 0.5200 939.8500 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 935.7500 0.5200 935.8500 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 931.7500 0.5200 931.8500 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 927.7500 0.5200 927.8500 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 923.7500 0.5200 923.8500 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 919.7500 0.5200 919.8500 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 915.7500 0.5200 915.8500 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 911.7500 0.5200 911.8500 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 907.7500 0.5200 907.8500 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 903.7500 0.5200 903.8500 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 899.7500 0.5200 899.8500 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 895.7500 0.5200 895.8500 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 891.7500 0.5200 891.8500 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 887.7500 0.5200 887.8500 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 883.7500 0.5200 883.8500 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 879.7500 0.5200 879.8500 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 875.7500 0.5200 875.8500 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 871.7500 0.5200 871.8500 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 867.7500 0.5200 867.8500 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 863.7500 0.5200 863.8500 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 859.7500 0.5200 859.8500 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 855.7500 0.5200 855.8500 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 851.7500 0.5200 851.8500 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 847.7500 0.5200 847.8500 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 843.7500 0.5200 843.8500 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 839.7500 0.5200 839.8500 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 835.7500 0.5200 835.8500 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 831.7500 0.5200 831.8500 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 827.7500 0.5200 827.8500 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 823.7500 0.5200 823.8500 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 819.7500 0.5200 819.8500 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 815.7500 0.5200 815.8500 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 811.7500 0.5200 811.8500 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 807.7500 0.5200 807.8500 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 803.7500 0.5200 803.8500 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 799.7500 0.5200 799.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 795.7500 0.5200 795.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 791.7500 0.5200 791.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 787.7500 0.5200 787.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 783.7500 0.5200 783.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 779.7500 0.5200 779.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 775.7500 0.5200 775.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 771.7500 0.5200 771.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 767.7500 0.5200 767.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 763.7500 0.5200 763.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 759.7500 0.5200 759.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 755.7500 0.5200 755.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 751.7500 0.5200 751.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 747.7500 0.5200 747.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 743.7500 0.5200 743.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 739.7500 0.5200 739.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 735.7500 0.5200 735.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 731.7500 0.5200 731.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 727.7500 0.5200 727.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 723.7500 0.5200 723.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 719.7500 0.5200 719.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 715.7500 0.5200 715.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 711.7500 0.5200 711.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 707.7500 0.5200 707.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 703.7500 0.5200 703.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 699.7500 0.5200 699.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 695.7500 0.5200 695.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 691.7500 0.5200 691.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 687.7500 0.5200 687.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 683.7500 0.5200 683.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 679.7500 0.5200 679.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 675.7500 0.5200 675.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 671.7500 0.5200 671.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 667.7500 0.5200 667.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 663.7500 0.5200 663.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 659.7500 0.5200 659.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 655.7500 0.5200 655.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 651.7500 0.5200 651.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 647.7500 0.5200 647.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 643.7500 0.5200 643.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 639.7500 0.5200 639.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 635.7500 0.5200 635.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 631.7500 0.5200 631.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 627.7500 0.5200 627.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 623.7500 0.5200 623.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 619.7500 0.5200 619.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 615.7500 0.5200 615.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 611.7500 0.5200 611.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 607.7500 0.5200 607.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 603.7500 0.5200 603.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 599.7500 0.5200 599.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 595.7500 0.5200 595.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 591.7500 0.5200 591.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 587.7500 0.5200 587.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 583.7500 0.5200 583.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 579.7500 0.5200 579.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 575.7500 0.5200 575.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 571.7500 0.5200 571.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 567.7500 0.5200 567.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 563.7500 0.5200 563.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 559.7500 0.5200 559.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 555.7500 0.5200 555.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 551.7500 0.5200 551.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 547.7500 0.5200 547.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 444.1500 1020.0000 444.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 448.1500 1020.0000 448.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 452.1500 1020.0000 452.2500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 456.1500 1020.0000 456.2500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 460.1500 1020.0000 460.2500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 464.1500 1020.0000 464.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 468.1500 1020.0000 468.2500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 472.1500 1020.0000 472.2500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 476.1500 1020.0000 476.2500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 480.1500 1020.0000 480.2500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 484.1500 1020.0000 484.2500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 488.1500 1020.0000 488.2500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 492.1500 1020.0000 492.2500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 496.1500 1020.0000 496.2500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 500.1500 1020.0000 500.2500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 504.1500 1020.0000 504.2500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 508.1500 1020.0000 508.2500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 512.1500 1020.0000 512.2500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 516.1500 1020.0000 516.2500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 520.1500 1020.0000 520.2500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 524.1500 1020.0000 524.2500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 528.1500 1020.0000 528.2500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 532.1500 1020.0000 532.2500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 536.1500 1020.0000 536.2500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 540.1500 1020.0000 540.2500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 544.1500 1020.0000 544.2500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 548.1500 1020.0000 548.2500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 552.1500 1020.0000 552.2500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 556.1500 1020.0000 556.2500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 560.1500 1020.0000 560.2500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 564.1500 1020.0000 564.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 568.1500 1020.0000 568.2500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 572.1500 1020.0000 572.2500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 576.1500 1020.0000 576.2500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 580.1500 1020.0000 580.2500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 584.1500 1020.0000 584.2500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 588.1500 1020.0000 588.2500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 592.1500 1020.0000 592.2500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 596.1500 1020.0000 596.2500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 600.1500 1020.0000 600.2500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 604.1500 1020.0000 604.2500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 608.1500 1020.0000 608.2500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 612.1500 1020.0000 612.2500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 616.1500 1020.0000 616.2500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 620.1500 1020.0000 620.2500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 624.1500 1020.0000 624.2500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 628.1500 1020.0000 628.2500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 632.1500 1020.0000 632.2500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 636.1500 1020.0000 636.2500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 640.1500 1020.0000 640.2500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 644.1500 1020.0000 644.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 648.1500 1020.0000 648.2500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 652.1500 1020.0000 652.2500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 656.1500 1020.0000 656.2500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 660.1500 1020.0000 660.2500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 664.1500 1020.0000 664.2500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 668.1500 1020.0000 668.2500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 672.1500 1020.0000 672.2500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 676.1500 1020.0000 676.2500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 680.1500 1020.0000 680.2500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 684.1500 1020.0000 684.2500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 688.1500 1020.0000 688.2500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 692.1500 1020.0000 692.2500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 696.1500 1020.0000 696.2500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 700.1500 1020.0000 700.2500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 704.1500 1020.0000 704.2500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 708.1500 1020.0000 708.2500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 712.1500 1020.0000 712.2500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 716.1500 1020.0000 716.2500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 720.1500 1020.0000 720.2500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 724.1500 1020.0000 724.2500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 728.1500 1020.0000 728.2500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 732.1500 1020.0000 732.2500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 736.1500 1020.0000 736.2500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 740.1500 1020.0000 740.2500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 744.1500 1020.0000 744.2500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 748.1500 1020.0000 748.2500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 752.1500 1020.0000 752.2500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 756.1500 1020.0000 756.2500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 760.1500 1020.0000 760.2500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 764.1500 1020.0000 764.2500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 768.1500 1020.0000 768.2500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 772.1500 1020.0000 772.2500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 776.1500 1020.0000 776.2500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 780.1500 1020.0000 780.2500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 784.1500 1020.0000 784.2500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 788.1500 1020.0000 788.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 792.1500 1020.0000 792.2500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 796.1500 1020.0000 796.2500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 800.1500 1020.0000 800.2500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 804.1500 1020.0000 804.2500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 808.1500 1020.0000 808.2500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 812.1500 1020.0000 812.2500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 816.1500 1020.0000 816.2500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 820.1500 1020.0000 820.2500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 824.1500 1020.0000 824.2500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 828.1500 1020.0000 828.2500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 832.1500 1020.0000 832.2500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 836.1500 1020.0000 836.2500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 840.1500 1020.0000 840.2500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 844.1500 1020.0000 844.2500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 848.1500 1020.0000 848.2500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 852.1500 1020.0000 852.2500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 856.1500 1020.0000 856.2500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 860.1500 1020.0000 860.2500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 864.1500 1020.0000 864.2500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 868.1500 1020.0000 868.2500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 872.1500 1020.0000 872.2500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 876.1500 1020.0000 876.2500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 880.1500 1020.0000 880.2500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 884.1500 1020.0000 884.2500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 888.1500 1020.0000 888.2500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 892.1500 1020.0000 892.2500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 896.1500 1020.0000 896.2500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 900.1500 1020.0000 900.2500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 904.1500 1020.0000 904.2500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 908.1500 1020.0000 908.2500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 912.1500 1020.0000 912.2500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 916.1500 1020.0000 916.2500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 920.1500 1020.0000 920.2500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 924.1500 1020.0000 924.2500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 928.1500 1020.0000 928.2500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 932.1500 1020.0000 932.2500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 936.1500 1020.0000 936.2500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 940.1500 1020.0000 940.2500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 944.1500 1020.0000 944.2500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 948.1500 1020.0000 948.2500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 952.1500 1020.0000 952.2500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 956.1500 1020.0000 956.2500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 960.1500 1020.0000 960.2500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 964.1500 1020.0000 964.2500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 968.1500 1020.0000 968.2500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 972.1500 1020.0000 972.2500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 976.1500 1020.0000 976.2500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 980.1500 1020.0000 980.2500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 984.1500 1020.0000 984.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 988.1500 1020.0000 988.2500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 992.1500 1020.0000 992.2500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 996.1500 1020.0000 996.2500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1000.1500 1020.0000 1000.2500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1004.1500 1020.0000 1004.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1008.1500 1020.0000 1008.2500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1012.1500 1020.0000 1012.2500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1016.1500 1020.0000 1016.2500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1020.1500 1020.0000 1020.2500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1024.1500 1020.0000 1024.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1028.1500 1020.0000 1028.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1032.1500 1020.0000 1032.2500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1036.1500 1020.0000 1036.2500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1040.1500 1020.0000 1040.2500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1044.1500 1020.0000 1044.2500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1048.1500 1020.0000 1048.2500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1052.1500 1020.0000 1052.2500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1056.1500 1020.0000 1056.2500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1060.1500 1020.0000 1060.2500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1064.1500 1020.0000 1064.2500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1068.1500 1020.0000 1068.2500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1072.1500 1020.0000 1072.2500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1076.1500 1020.0000 1076.2500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1019.4800 1080.1500 1020.0000 1080.2500 ;
    END
  END out[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 543.7500 0.5200 543.8500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 539.7500 0.5200 539.8500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 535.7500 0.5200 535.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 531.7500 0.5200 531.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 527.7500 0.5200 527.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 523.7500 0.5200 523.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 519.7500 0.5200 519.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 515.7500 0.5200 515.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 511.7500 0.5200 511.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 507.7500 0.5200 507.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 503.7500 0.5200 503.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 499.7500 0.5200 499.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 495.7500 0.5200 495.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 491.7500 0.5200 491.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 487.7500 0.5200 487.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 483.7500 0.5200 483.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 479.7500 0.5200 479.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 475.7500 0.5200 475.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 471.7500 0.5200 471.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 1059.7500 0.5200 1059.8500 ;
    END
  END reset
  PIN fifo_ext_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 467.7500 0.5200 467.8500 ;
    END
  END fifo_ext_rd
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 1000.0000 10.0000 1002.0000 1610.0000 ;
        RECT 890.0000 10.0000 892.0000 1610.0000 ;
        RECT 780.0000 10.0000 782.0000 1610.0000 ;
        RECT 670.0000 10.0000 672.0000 1610.0000 ;
        RECT 560.0000 10.0000 562.0000 1610.0000 ;
        RECT 450.0000 10.0000 452.0000 1610.0000 ;
        RECT 340.0000 10.0000 342.0000 1610.0000 ;
        RECT 230.0000 10.0000 232.0000 1610.0000 ;
        RECT 120.0000 10.0000 122.0000 1610.0000 ;
        RECT 10.0000 10.0000 12.0000 1610.0000 ;
        RECT 99.3850 202.4350 99.7150 202.7650 ;
        RECT 99.3850 101.6350 99.7150 101.9650 ;
        RECT 99.3850 105.2350 99.7150 105.5650 ;
        RECT 99.3850 108.8350 99.7150 109.1650 ;
        RECT 99.3850 112.4350 99.7150 112.7650 ;
        RECT 99.3850 116.0350 99.7150 116.3650 ;
        RECT 99.3850 119.6350 99.7150 119.9650 ;
        RECT 99.3850 123.2350 99.7150 123.5650 ;
        RECT 99.3850 126.8350 99.7150 127.1650 ;
        RECT 99.3850 130.4350 99.7150 130.7650 ;
        RECT 99.3850 134.0350 99.7150 134.3650 ;
        RECT 99.3850 137.6350 99.7150 137.9650 ;
        RECT 99.3850 141.2350 99.7150 141.5650 ;
        RECT 99.3850 144.8350 99.7150 145.1650 ;
        RECT 99.3850 148.4350 99.7150 148.7650 ;
        RECT 99.3850 152.0350 99.7150 152.3650 ;
        RECT 99.3850 155.6350 99.7150 155.9650 ;
        RECT 99.3850 159.2350 99.7150 159.5650 ;
        RECT 99.3850 162.8350 99.7150 163.1650 ;
        RECT 99.3850 166.4350 99.7150 166.7650 ;
        RECT 99.3850 170.0350 99.7150 170.3650 ;
        RECT 99.3850 173.6350 99.7150 173.9650 ;
        RECT 99.3850 177.2350 99.7150 177.5650 ;
        RECT 99.3850 180.8350 99.7150 181.1650 ;
        RECT 99.3850 184.4350 99.7150 184.7650 ;
        RECT 99.3850 188.0350 99.7150 188.3650 ;
        RECT 99.3850 195.2350 99.7150 195.5650 ;
        RECT 99.3850 191.6350 99.7150 191.9650 ;
        RECT 99.3850 198.8350 99.7150 199.1650 ;
        RECT 99.3850 252.8350 99.7150 253.1650 ;
        RECT 99.3850 227.6350 99.7150 227.9650 ;
        RECT 99.3850 206.0350 99.7150 206.3650 ;
        RECT 99.3850 209.6350 99.7150 209.9650 ;
        RECT 99.3850 213.2350 99.7150 213.5650 ;
        RECT 99.3850 220.4350 99.7150 220.7650 ;
        RECT 99.3850 216.8350 99.7150 217.1650 ;
        RECT 99.3850 224.0350 99.7150 224.3650 ;
        RECT 99.3850 231.2350 99.7150 231.5650 ;
        RECT 99.3850 234.8350 99.7150 235.1650 ;
        RECT 99.3850 238.4350 99.7150 238.7650 ;
        RECT 99.3850 245.6350 99.7150 245.9650 ;
        RECT 99.3850 242.0350 99.7150 242.3650 ;
        RECT 99.3850 249.2350 99.7150 249.5650 ;
        RECT 99.3850 256.4350 99.7150 256.7650 ;
        RECT 99.3850 260.0350 99.7150 260.3650 ;
        RECT 99.3850 263.6350 99.7150 263.9650 ;
        RECT 99.3850 267.2350 99.7150 267.5650 ;
        RECT 99.3850 270.8350 99.7150 271.1650 ;
        RECT 99.3850 274.4350 99.7150 274.7650 ;
        RECT 99.3850 278.0350 99.7150 278.3650 ;
        RECT 99.3850 281.6350 99.7150 281.9650 ;
        RECT 99.3850 285.2350 99.7150 285.5650 ;
        RECT 99.3850 288.8350 99.7150 289.1650 ;
        RECT 99.3850 292.4350 99.7150 292.7650 ;
        RECT 99.3850 296.0350 99.7150 296.3650 ;
        RECT 99.3850 299.6350 99.7150 299.9650 ;
        RECT 99.3850 303.2350 99.7150 303.5650 ;
        RECT 99.3850 306.8350 99.7150 307.1650 ;
        RECT 99.3850 310.4350 99.7150 310.7650 ;
        RECT 99.3850 314.0350 99.7150 314.3650 ;
        RECT 99.3850 317.6350 99.7150 317.9650 ;
        RECT 99.3850 321.2350 99.7150 321.5650 ;
        RECT 99.3850 324.8350 99.7150 325.1650 ;
        RECT 99.3850 328.4350 99.7150 328.7650 ;
        RECT 99.3850 332.0350 99.7150 332.3650 ;
        RECT 99.3850 335.6350 99.7150 335.9650 ;
        RECT 99.3850 339.2350 99.7150 339.5650 ;
        RECT 99.3850 342.8350 99.7150 343.1650 ;
        RECT 99.3850 346.4350 99.7150 346.7650 ;
        RECT 99.3850 350.0350 99.7150 350.3650 ;
        RECT 99.3850 353.6350 99.7150 353.9650 ;
        RECT 99.3850 357.2350 99.7150 357.5650 ;
        RECT 99.3850 360.8350 99.7150 361.1650 ;
        RECT 99.3850 364.4350 99.7150 364.7650 ;
        RECT 99.3850 368.0350 99.7150 368.3650 ;
        RECT 99.3850 371.6350 99.7150 371.9650 ;
        RECT 99.3850 375.2350 99.7150 375.5650 ;
        RECT 99.3850 378.8350 99.7150 379.1650 ;
        RECT 99.3850 382.4350 99.7150 382.7650 ;
        RECT 99.3850 386.0350 99.7150 386.3650 ;
        RECT 99.3850 389.6350 99.7150 389.9650 ;
        RECT 99.3850 393.2350 99.7150 393.5650 ;
        RECT 99.3850 396.8350 99.7150 397.1650 ;
        RECT 99.3850 400.4350 99.7150 400.7650 ;
        RECT 99.3850 404.0350 99.7150 404.3650 ;
        RECT 99.3850 411.2350 99.7150 411.5650 ;
        RECT 99.3850 407.6350 99.7150 407.9650 ;
        RECT 99.3850 414.8350 99.7150 415.1650 ;
        RECT 99.3850 418.4350 99.7150 418.7650 ;
        RECT 99.3850 422.0350 99.7150 422.3650 ;
        RECT 99.3850 425.6350 99.7150 425.9650 ;
        RECT 99.3850 429.2350 99.7150 429.5650 ;
        RECT 99.3850 436.4350 99.7150 436.7650 ;
        RECT 99.3850 432.8350 99.7150 433.1650 ;
        RECT 99.3850 440.0350 99.7150 440.3650 ;
        RECT 99.3850 443.6350 99.7150 443.9650 ;
        RECT 99.3850 447.2350 99.7150 447.5650 ;
        RECT 99.3850 450.8350 99.7150 451.1650 ;
        RECT 99.3850 454.4350 99.7150 454.7650 ;
        RECT 99.3850 461.6350 99.7150 461.9650 ;
        RECT 99.3850 458.0350 99.7150 458.3650 ;
        RECT 99.3850 465.2350 99.7150 465.5650 ;
        RECT 99.3850 468.8350 99.7150 469.1650 ;
        RECT 99.3850 472.4350 99.7150 472.7650 ;
        RECT 99.3850 476.0350 99.7150 476.3650 ;
        RECT 99.3850 479.6350 99.7150 479.9650 ;
        RECT 99.3850 483.2350 99.7150 483.5650 ;
        RECT 99.3850 486.8350 99.7150 487.1650 ;
        RECT 99.3850 490.4350 99.7150 490.7650 ;
        RECT 99.3850 494.0350 99.7150 494.3650 ;
        RECT 99.3850 497.6350 99.7150 497.9650 ;
        RECT 99.3850 501.2350 99.7150 501.5650 ;
        RECT 99.3850 504.8350 99.7150 505.1650 ;
        RECT 99.3850 508.4350 99.7150 508.7650 ;
        RECT 99.3850 512.0350 99.7150 512.3650 ;
        RECT 99.3850 515.6350 99.7150 515.9650 ;
        RECT 99.3850 519.2350 99.7150 519.5650 ;
        RECT 99.3850 602.0350 99.7150 602.3650 ;
        RECT 99.3850 605.6350 99.7150 605.9650 ;
        RECT 99.3850 620.0350 99.7150 620.3650 ;
        RECT 99.3850 612.8350 99.7150 613.1650 ;
        RECT 99.3850 609.2350 99.7150 609.5650 ;
        RECT 99.3850 616.4350 99.7150 616.7650 ;
        RECT 99.3850 623.6350 99.7150 623.9650 ;
        RECT 99.3850 627.2350 99.7150 627.5650 ;
        RECT 99.3850 630.8350 99.7150 631.1650 ;
        RECT 99.3850 645.2350 99.7150 645.5650 ;
        RECT 99.3850 638.0350 99.7150 638.3650 ;
        RECT 99.3850 634.4350 99.7150 634.7650 ;
        RECT 99.3850 641.6350 99.7150 641.9650 ;
        RECT 99.3850 648.8350 99.7150 649.1650 ;
        RECT 99.3850 652.4350 99.7150 652.7650 ;
        RECT 99.3850 656.0350 99.7150 656.3650 ;
        RECT 99.3850 659.6350 99.7150 659.9650 ;
        RECT 99.3850 663.2350 99.7150 663.5650 ;
        RECT 99.3850 666.8350 99.7150 667.1650 ;
        RECT 99.3850 670.4350 99.7150 670.7650 ;
        RECT 99.3850 674.0350 99.7150 674.3650 ;
        RECT 99.3850 677.6350 99.7150 677.9650 ;
        RECT 99.3850 681.2350 99.7150 681.5650 ;
        RECT 99.3850 684.8350 99.7150 685.1650 ;
        RECT 99.3850 688.4350 99.7150 688.7650 ;
        RECT 99.3850 692.0350 99.7150 692.3650 ;
        RECT 99.3850 695.6350 99.7150 695.9650 ;
        RECT 99.3850 699.2350 99.7150 699.5650 ;
        RECT 99.3850 702.8350 99.7150 703.1650 ;
        RECT 99.3850 706.4350 99.7150 706.7650 ;
        RECT 99.3850 710.0350 99.7150 710.3650 ;
        RECT 99.3850 713.6350 99.7150 713.9650 ;
        RECT 99.3850 717.2350 99.7150 717.5650 ;
        RECT 99.3850 720.8350 99.7150 721.1650 ;
        RECT 99.3850 724.4350 99.7150 724.7650 ;
        RECT 99.3850 728.0350 99.7150 728.3650 ;
        RECT 99.3850 731.6350 99.7150 731.9650 ;
        RECT 99.3850 735.2350 99.7150 735.5650 ;
        RECT 99.3850 738.8350 99.7150 739.1650 ;
        RECT 99.3850 742.4350 99.7150 742.7650 ;
        RECT 99.3850 746.0350 99.7150 746.3650 ;
        RECT 99.3850 749.6350 99.7150 749.9650 ;
        RECT 99.3850 753.2350 99.7150 753.5650 ;
        RECT 99.3850 756.8350 99.7150 757.1650 ;
        RECT 99.3850 760.4350 99.7150 760.7650 ;
        RECT 99.3850 764.0350 99.7150 764.3650 ;
        RECT 99.3850 767.6350 99.7150 767.9650 ;
        RECT 99.3850 771.2350 99.7150 771.5650 ;
        RECT 99.3850 774.8350 99.7150 775.1650 ;
        RECT 99.3850 778.4350 99.7150 778.7650 ;
        RECT 99.3850 782.0350 99.7150 782.3650 ;
        RECT 99.3850 785.6350 99.7150 785.9650 ;
        RECT 99.3850 789.2350 99.7150 789.5650 ;
        RECT 99.3850 792.8350 99.7150 793.1650 ;
        RECT 99.3850 796.4350 99.7150 796.7650 ;
        RECT 99.3850 803.6350 99.7150 803.9650 ;
        RECT 99.3850 800.0350 99.7150 800.3650 ;
        RECT 99.3850 807.2350 99.7150 807.5650 ;
        RECT 920.1200 202.4350 920.4500 202.7650 ;
        RECT 920.1200 101.6350 920.4500 101.9650 ;
        RECT 920.1200 105.2350 920.4500 105.5650 ;
        RECT 920.1200 108.8350 920.4500 109.1650 ;
        RECT 920.1200 112.4350 920.4500 112.7650 ;
        RECT 920.1200 116.0350 920.4500 116.3650 ;
        RECT 920.1200 119.6350 920.4500 119.9650 ;
        RECT 920.1200 123.2350 920.4500 123.5650 ;
        RECT 920.1200 126.8350 920.4500 127.1650 ;
        RECT 920.1200 130.4350 920.4500 130.7650 ;
        RECT 920.1200 134.0350 920.4500 134.3650 ;
        RECT 920.1200 137.6350 920.4500 137.9650 ;
        RECT 920.1200 141.2350 920.4500 141.5650 ;
        RECT 920.1200 144.8350 920.4500 145.1650 ;
        RECT 920.1200 148.4350 920.4500 148.7650 ;
        RECT 920.1200 152.0350 920.4500 152.3650 ;
        RECT 920.1200 155.6350 920.4500 155.9650 ;
        RECT 920.1200 159.2350 920.4500 159.5650 ;
        RECT 920.1200 162.8350 920.4500 163.1650 ;
        RECT 920.1200 166.4350 920.4500 166.7650 ;
        RECT 920.1200 170.0350 920.4500 170.3650 ;
        RECT 920.1200 173.6350 920.4500 173.9650 ;
        RECT 920.1200 177.2350 920.4500 177.5650 ;
        RECT 920.1200 180.8350 920.4500 181.1650 ;
        RECT 920.1200 184.4350 920.4500 184.7650 ;
        RECT 920.1200 188.0350 920.4500 188.3650 ;
        RECT 920.1200 195.2350 920.4500 195.5650 ;
        RECT 920.1200 191.6350 920.4500 191.9650 ;
        RECT 920.1200 198.8350 920.4500 199.1650 ;
        RECT 920.1200 252.8350 920.4500 253.1650 ;
        RECT 920.1200 227.6350 920.4500 227.9650 ;
        RECT 920.1200 206.0350 920.4500 206.3650 ;
        RECT 920.1200 209.6350 920.4500 209.9650 ;
        RECT 920.1200 213.2350 920.4500 213.5650 ;
        RECT 920.1200 220.4350 920.4500 220.7650 ;
        RECT 920.1200 216.8350 920.4500 217.1650 ;
        RECT 920.1200 224.0350 920.4500 224.3650 ;
        RECT 920.1200 231.2350 920.4500 231.5650 ;
        RECT 920.1200 234.8350 920.4500 235.1650 ;
        RECT 920.1200 238.4350 920.4500 238.7650 ;
        RECT 920.1200 245.6350 920.4500 245.9650 ;
        RECT 920.1200 242.0350 920.4500 242.3650 ;
        RECT 920.1200 249.2350 920.4500 249.5650 ;
        RECT 920.1200 256.4350 920.4500 256.7650 ;
        RECT 920.1200 260.0350 920.4500 260.3650 ;
        RECT 920.1200 263.6350 920.4500 263.9650 ;
        RECT 920.1200 267.2350 920.4500 267.5650 ;
        RECT 920.1200 270.8350 920.4500 271.1650 ;
        RECT 920.1200 274.4350 920.4500 274.7650 ;
        RECT 920.1200 278.0350 920.4500 278.3650 ;
        RECT 920.1200 281.6350 920.4500 281.9650 ;
        RECT 920.1200 285.2350 920.4500 285.5650 ;
        RECT 920.1200 288.8350 920.4500 289.1650 ;
        RECT 920.1200 292.4350 920.4500 292.7650 ;
        RECT 920.1200 296.0350 920.4500 296.3650 ;
        RECT 920.1200 299.6350 920.4500 299.9650 ;
        RECT 920.1200 303.2350 920.4500 303.5650 ;
        RECT 920.1200 306.8350 920.4500 307.1650 ;
        RECT 920.1200 310.4350 920.4500 310.7650 ;
        RECT 920.1200 314.0350 920.4500 314.3650 ;
        RECT 920.1200 317.6350 920.4500 317.9650 ;
        RECT 920.1200 321.2350 920.4500 321.5650 ;
        RECT 920.1200 324.8350 920.4500 325.1650 ;
        RECT 920.1200 328.4350 920.4500 328.7650 ;
        RECT 920.1200 332.0350 920.4500 332.3650 ;
        RECT 920.1200 335.6350 920.4500 335.9650 ;
        RECT 920.1200 339.2350 920.4500 339.5650 ;
        RECT 920.1200 342.8350 920.4500 343.1650 ;
        RECT 920.1200 346.4350 920.4500 346.7650 ;
        RECT 920.1200 350.0350 920.4500 350.3650 ;
        RECT 920.1200 353.6350 920.4500 353.9650 ;
        RECT 920.1200 357.2350 920.4500 357.5650 ;
        RECT 920.1200 360.8350 920.4500 361.1650 ;
        RECT 920.1200 364.4350 920.4500 364.7650 ;
        RECT 920.1200 368.0350 920.4500 368.3650 ;
        RECT 920.1200 371.6350 920.4500 371.9650 ;
        RECT 920.1200 375.2350 920.4500 375.5650 ;
        RECT 920.1200 378.8350 920.4500 379.1650 ;
        RECT 920.1200 382.4350 920.4500 382.7650 ;
        RECT 920.1200 386.0350 920.4500 386.3650 ;
        RECT 920.1200 389.6350 920.4500 389.9650 ;
        RECT 920.1200 393.2350 920.4500 393.5650 ;
        RECT 920.1200 396.8350 920.4500 397.1650 ;
        RECT 920.1200 400.4350 920.4500 400.7650 ;
        RECT 920.1200 404.0350 920.4500 404.3650 ;
        RECT 920.1200 411.2350 920.4500 411.5650 ;
        RECT 920.1200 407.6350 920.4500 407.9650 ;
        RECT 920.1200 414.8350 920.4500 415.1650 ;
        RECT 920.1200 418.4350 920.4500 418.7650 ;
        RECT 920.1200 422.0350 920.4500 422.3650 ;
        RECT 920.1200 425.6350 920.4500 425.9650 ;
        RECT 920.1200 429.2350 920.4500 429.5650 ;
        RECT 920.1200 436.4350 920.4500 436.7650 ;
        RECT 920.1200 432.8350 920.4500 433.1650 ;
        RECT 920.1200 440.0350 920.4500 440.3650 ;
        RECT 920.1200 443.6350 920.4500 443.9650 ;
        RECT 920.1200 447.2350 920.4500 447.5650 ;
        RECT 920.1200 450.8350 920.4500 451.1650 ;
        RECT 920.1200 454.4350 920.4500 454.7650 ;
        RECT 920.1200 461.6350 920.4500 461.9650 ;
        RECT 920.1200 458.0350 920.4500 458.3650 ;
        RECT 920.1200 465.2350 920.4500 465.5650 ;
        RECT 920.1200 468.8350 920.4500 469.1650 ;
        RECT 920.1200 472.4350 920.4500 472.7650 ;
        RECT 920.1200 476.0350 920.4500 476.3650 ;
        RECT 920.1200 479.6350 920.4500 479.9650 ;
        RECT 920.1200 483.2350 920.4500 483.5650 ;
        RECT 920.1200 486.8350 920.4500 487.1650 ;
        RECT 920.1200 490.4350 920.4500 490.7650 ;
        RECT 920.1200 494.0350 920.4500 494.3650 ;
        RECT 920.1200 497.6350 920.4500 497.9650 ;
        RECT 920.1200 501.2350 920.4500 501.5650 ;
        RECT 920.1200 504.8350 920.4500 505.1650 ;
        RECT 920.1200 508.4350 920.4500 508.7650 ;
        RECT 920.1200 512.0350 920.4500 512.3650 ;
        RECT 920.1200 515.6350 920.4500 515.9650 ;
        RECT 920.1200 519.2350 920.4500 519.5650 ;
        RECT 920.1200 602.0350 920.4500 602.3650 ;
        RECT 920.1200 605.6350 920.4500 605.9650 ;
        RECT 920.1200 620.0350 920.4500 620.3650 ;
        RECT 920.1200 612.8350 920.4500 613.1650 ;
        RECT 920.1200 609.2350 920.4500 609.5650 ;
        RECT 920.1200 616.4350 920.4500 616.7650 ;
        RECT 920.1200 623.6350 920.4500 623.9650 ;
        RECT 920.1200 627.2350 920.4500 627.5650 ;
        RECT 920.1200 630.8350 920.4500 631.1650 ;
        RECT 920.1200 645.2350 920.4500 645.5650 ;
        RECT 920.1200 638.0350 920.4500 638.3650 ;
        RECT 920.1200 634.4350 920.4500 634.7650 ;
        RECT 920.1200 641.6350 920.4500 641.9650 ;
        RECT 920.1200 648.8350 920.4500 649.1650 ;
        RECT 920.1200 652.4350 920.4500 652.7650 ;
        RECT 920.1200 656.0350 920.4500 656.3650 ;
        RECT 920.1200 659.6350 920.4500 659.9650 ;
        RECT 920.1200 663.2350 920.4500 663.5650 ;
        RECT 920.1200 666.8350 920.4500 667.1650 ;
        RECT 920.1200 670.4350 920.4500 670.7650 ;
        RECT 920.1200 674.0350 920.4500 674.3650 ;
        RECT 920.1200 677.6350 920.4500 677.9650 ;
        RECT 920.1200 681.2350 920.4500 681.5650 ;
        RECT 920.1200 684.8350 920.4500 685.1650 ;
        RECT 920.1200 688.4350 920.4500 688.7650 ;
        RECT 920.1200 692.0350 920.4500 692.3650 ;
        RECT 920.1200 695.6350 920.4500 695.9650 ;
        RECT 920.1200 699.2350 920.4500 699.5650 ;
        RECT 920.1200 702.8350 920.4500 703.1650 ;
        RECT 920.1200 706.4350 920.4500 706.7650 ;
        RECT 920.1200 710.0350 920.4500 710.3650 ;
        RECT 920.1200 713.6350 920.4500 713.9650 ;
        RECT 920.1200 717.2350 920.4500 717.5650 ;
        RECT 920.1200 720.8350 920.4500 721.1650 ;
        RECT 920.1200 724.4350 920.4500 724.7650 ;
        RECT 920.1200 728.0350 920.4500 728.3650 ;
        RECT 920.1200 731.6350 920.4500 731.9650 ;
        RECT 920.1200 735.2350 920.4500 735.5650 ;
        RECT 920.1200 738.8350 920.4500 739.1650 ;
        RECT 920.1200 742.4350 920.4500 742.7650 ;
        RECT 920.1200 746.0350 920.4500 746.3650 ;
        RECT 920.1200 749.6350 920.4500 749.9650 ;
        RECT 920.1200 753.2350 920.4500 753.5650 ;
        RECT 920.1200 756.8350 920.4500 757.1650 ;
        RECT 920.1200 760.4350 920.4500 760.7650 ;
        RECT 920.1200 764.0350 920.4500 764.3650 ;
        RECT 920.1200 767.6350 920.4500 767.9650 ;
        RECT 920.1200 771.2350 920.4500 771.5650 ;
        RECT 920.1200 774.8350 920.4500 775.1650 ;
        RECT 920.1200 778.4350 920.4500 778.7650 ;
        RECT 920.1200 782.0350 920.4500 782.3650 ;
        RECT 920.1200 785.6350 920.4500 785.9650 ;
        RECT 920.1200 789.2350 920.4500 789.5650 ;
        RECT 920.1200 792.8350 920.4500 793.1650 ;
        RECT 920.1200 796.4350 920.4500 796.7650 ;
        RECT 920.1200 803.6350 920.4500 803.9650 ;
        RECT 920.1200 800.0350 920.4500 800.3650 ;
        RECT 920.1200 807.2350 920.4500 807.5650 ;
        RECT 99.3850 1012.4350 99.7150 1012.7650 ;
        RECT 99.3850 810.8350 99.7150 811.1650 ;
        RECT 99.3850 814.4350 99.7150 814.7650 ;
        RECT 99.3850 818.0350 99.7150 818.3650 ;
        RECT 99.3850 821.6350 99.7150 821.9650 ;
        RECT 99.3850 828.8350 99.7150 829.1650 ;
        RECT 99.3850 825.2350 99.7150 825.5650 ;
        RECT 99.3850 832.4350 99.7150 832.7650 ;
        RECT 99.3850 836.0350 99.7150 836.3650 ;
        RECT 99.3850 839.6350 99.7150 839.9650 ;
        RECT 99.3850 843.2350 99.7150 843.5650 ;
        RECT 99.3850 846.8350 99.7150 847.1650 ;
        RECT 99.3850 854.0350 99.7150 854.3650 ;
        RECT 99.3850 850.4350 99.7150 850.7650 ;
        RECT 99.3850 857.6350 99.7150 857.9650 ;
        RECT 99.3850 861.2350 99.7150 861.5650 ;
        RECT 99.3850 864.8350 99.7150 865.1650 ;
        RECT 99.3850 868.4350 99.7150 868.7650 ;
        RECT 99.3850 872.0350 99.7150 872.3650 ;
        RECT 99.3850 875.6350 99.7150 875.9650 ;
        RECT 99.3850 879.2350 99.7150 879.5650 ;
        RECT 99.3850 882.8350 99.7150 883.1650 ;
        RECT 99.3850 886.4350 99.7150 886.7650 ;
        RECT 99.3850 890.0350 99.7150 890.3650 ;
        RECT 99.3850 893.6350 99.7150 893.9650 ;
        RECT 99.3850 897.2350 99.7150 897.5650 ;
        RECT 99.3850 900.8350 99.7150 901.1650 ;
        RECT 99.3850 904.4350 99.7150 904.7650 ;
        RECT 99.3850 908.0350 99.7150 908.3650 ;
        RECT 99.3850 911.6350 99.7150 911.9650 ;
        RECT 99.3850 915.2350 99.7150 915.5650 ;
        RECT 99.3850 918.8350 99.7150 919.1650 ;
        RECT 99.3850 922.4350 99.7150 922.7650 ;
        RECT 99.3850 926.0350 99.7150 926.3650 ;
        RECT 99.3850 929.6350 99.7150 929.9650 ;
        RECT 99.3850 933.2350 99.7150 933.5650 ;
        RECT 99.3850 936.8350 99.7150 937.1650 ;
        RECT 99.3850 940.4350 99.7150 940.7650 ;
        RECT 99.3850 944.0350 99.7150 944.3650 ;
        RECT 99.3850 947.6350 99.7150 947.9650 ;
        RECT 99.3850 951.2350 99.7150 951.5650 ;
        RECT 99.3850 954.8350 99.7150 955.1650 ;
        RECT 99.3850 958.4350 99.7150 958.7650 ;
        RECT 99.3850 962.0350 99.7150 962.3650 ;
        RECT 99.3850 965.6350 99.7150 965.9650 ;
        RECT 99.3850 969.2350 99.7150 969.5650 ;
        RECT 99.3850 972.8350 99.7150 973.1650 ;
        RECT 99.3850 976.4350 99.7150 976.7650 ;
        RECT 99.3850 980.0350 99.7150 980.3650 ;
        RECT 99.3850 983.6350 99.7150 983.9650 ;
        RECT 99.3850 987.2350 99.7150 987.5650 ;
        RECT 99.3850 990.8350 99.7150 991.1650 ;
        RECT 99.3850 994.4350 99.7150 994.7650 ;
        RECT 99.3850 998.0350 99.7150 998.3650 ;
        RECT 99.3850 1005.2350 99.7150 1005.5650 ;
        RECT 99.3850 1001.6350 99.7150 1001.9650 ;
        RECT 99.3850 1008.8350 99.7150 1009.1650 ;
        RECT 99.3850 1016.0350 99.7150 1016.3650 ;
        RECT 99.3850 1019.6350 99.7150 1019.9650 ;
        RECT 99.3850 1102.4350 99.7150 1102.7650 ;
        RECT 99.3850 1106.0350 99.7150 1106.3650 ;
        RECT 99.3850 1109.6350 99.7150 1109.9650 ;
        RECT 99.3850 1113.2350 99.7150 1113.5650 ;
        RECT 99.3850 1116.8350 99.7150 1117.1650 ;
        RECT 99.3850 1120.4350 99.7150 1120.7650 ;
        RECT 99.3850 1124.0350 99.7150 1124.3650 ;
        RECT 99.3850 1127.6350 99.7150 1127.9650 ;
        RECT 99.3850 1131.2350 99.7150 1131.5650 ;
        RECT 99.3850 1134.8350 99.7150 1135.1650 ;
        RECT 99.3850 1138.4350 99.7150 1138.7650 ;
        RECT 99.3850 1142.0350 99.7150 1142.3650 ;
        RECT 99.3850 1145.6350 99.7150 1145.9650 ;
        RECT 99.3850 1149.2350 99.7150 1149.5650 ;
        RECT 99.3850 1152.8350 99.7150 1153.1650 ;
        RECT 99.3850 1156.4350 99.7150 1156.7650 ;
        RECT 99.3850 1160.0350 99.7150 1160.3650 ;
        RECT 99.3850 1163.6350 99.7150 1163.9650 ;
        RECT 99.3850 1167.2350 99.7150 1167.5650 ;
        RECT 99.3850 1170.8350 99.7150 1171.1650 ;
        RECT 99.3850 1174.4350 99.7150 1174.7650 ;
        RECT 99.3850 1178.0350 99.7150 1178.3650 ;
        RECT 99.3850 1181.6350 99.7150 1181.9650 ;
        RECT 99.3850 1185.2350 99.7150 1185.5650 ;
        RECT 99.3850 1188.8350 99.7150 1189.1650 ;
        RECT 99.3850 1192.4350 99.7150 1192.7650 ;
        RECT 99.3850 1196.0350 99.7150 1196.3650 ;
        RECT 99.3850 1199.6350 99.7150 1199.9650 ;
        RECT 99.3850 1203.2350 99.7150 1203.5650 ;
        RECT 99.3850 1206.8350 99.7150 1207.1650 ;
        RECT 99.3850 1210.4350 99.7150 1210.7650 ;
        RECT 99.3850 1214.0350 99.7150 1214.3650 ;
        RECT 99.3850 1221.2350 99.7150 1221.5650 ;
        RECT 99.3850 1217.6350 99.7150 1217.9650 ;
        RECT 99.3850 1224.8350 99.7150 1225.1650 ;
        RECT 99.3850 1228.4350 99.7150 1228.7650 ;
        RECT 99.3850 1232.0350 99.7150 1232.3650 ;
        RECT 99.3850 1235.6350 99.7150 1235.9650 ;
        RECT 99.3850 1239.2350 99.7150 1239.5650 ;
        RECT 99.3850 1246.4350 99.7150 1246.7650 ;
        RECT 99.3850 1242.8350 99.7150 1243.1650 ;
        RECT 99.3850 1250.0350 99.7150 1250.3650 ;
        RECT 99.3850 1253.6350 99.7150 1253.9650 ;
        RECT 99.3850 1257.2350 99.7150 1257.5650 ;
        RECT 99.3850 1260.8350 99.7150 1261.1650 ;
        RECT 99.3850 1264.4350 99.7150 1264.7650 ;
        RECT 99.3850 1271.6350 99.7150 1271.9650 ;
        RECT 99.3850 1268.0350 99.7150 1268.3650 ;
        RECT 99.3850 1275.2350 99.7150 1275.5650 ;
        RECT 99.3850 1278.8350 99.7150 1279.1650 ;
        RECT 99.3850 1282.4350 99.7150 1282.7650 ;
        RECT 99.3850 1286.0350 99.7150 1286.3650 ;
        RECT 99.3850 1289.6350 99.7150 1289.9650 ;
        RECT 99.3850 1293.2350 99.7150 1293.5650 ;
        RECT 99.3850 1296.8350 99.7150 1297.1650 ;
        RECT 99.3850 1300.4350 99.7150 1300.7650 ;
        RECT 99.3850 1304.0350 99.7150 1304.3650 ;
        RECT 99.3850 1307.6350 99.7150 1307.9650 ;
        RECT 99.3850 1311.2350 99.7150 1311.5650 ;
        RECT 99.3850 1314.8350 99.7150 1315.1650 ;
        RECT 99.3850 1318.4350 99.7150 1318.7650 ;
        RECT 99.3850 1322.0350 99.7150 1322.3650 ;
        RECT 99.3850 1325.6350 99.7150 1325.9650 ;
        RECT 99.3850 1329.2350 99.7150 1329.5650 ;
        RECT 99.3850 1332.8350 99.7150 1333.1650 ;
        RECT 99.3850 1336.4350 99.7150 1336.7650 ;
        RECT 99.3850 1340.0350 99.7150 1340.3650 ;
        RECT 99.3850 1343.6350 99.7150 1343.9650 ;
        RECT 99.3850 1347.2350 99.7150 1347.5650 ;
        RECT 99.3850 1350.8350 99.7150 1351.1650 ;
        RECT 99.3850 1354.4350 99.7150 1354.7650 ;
        RECT 99.3850 1358.0350 99.7150 1358.3650 ;
        RECT 99.3850 1361.6350 99.7150 1361.9650 ;
        RECT 99.3850 1365.2350 99.7150 1365.5650 ;
        RECT 99.3850 1368.8350 99.7150 1369.1650 ;
        RECT 99.3850 1372.4350 99.7150 1372.7650 ;
        RECT 99.3850 1376.0350 99.7150 1376.3650 ;
        RECT 99.3850 1379.6350 99.7150 1379.9650 ;
        RECT 99.3850 1383.2350 99.7150 1383.5650 ;
        RECT 99.3850 1386.8350 99.7150 1387.1650 ;
        RECT 99.3850 1390.4350 99.7150 1390.7650 ;
        RECT 99.3850 1404.8350 99.7150 1405.1650 ;
        RECT 99.3850 1394.0350 99.7150 1394.3650 ;
        RECT 99.3850 1397.6350 99.7150 1397.9650 ;
        RECT 99.3850 1401.2350 99.7150 1401.5650 ;
        RECT 99.3850 1408.4350 99.7150 1408.7650 ;
        RECT 99.3850 1412.0350 99.7150 1412.3650 ;
        RECT 99.3850 1415.6350 99.7150 1415.9650 ;
        RECT 99.3850 1430.0350 99.7150 1430.3650 ;
        RECT 99.3850 1422.8350 99.7150 1423.1650 ;
        RECT 99.3850 1419.2350 99.7150 1419.5650 ;
        RECT 99.3850 1426.4350 99.7150 1426.7650 ;
        RECT 99.3850 1433.6350 99.7150 1433.9650 ;
        RECT 99.3850 1437.2350 99.7150 1437.5650 ;
        RECT 99.3850 1440.8350 99.7150 1441.1650 ;
        RECT 99.3850 1455.2350 99.7150 1455.5650 ;
        RECT 99.3850 1448.0350 99.7150 1448.3650 ;
        RECT 99.3850 1444.4350 99.7150 1444.7650 ;
        RECT 99.3850 1451.6350 99.7150 1451.9650 ;
        RECT 99.3850 1458.8350 99.7150 1459.1650 ;
        RECT 99.3850 1462.4350 99.7150 1462.7650 ;
        RECT 99.3850 1466.0350 99.7150 1466.3650 ;
        RECT 99.3850 1469.6350 99.7150 1469.9650 ;
        RECT 99.3850 1473.2350 99.7150 1473.5650 ;
        RECT 99.3850 1476.8350 99.7150 1477.1650 ;
        RECT 99.3850 1480.4350 99.7150 1480.7650 ;
        RECT 99.3850 1484.0350 99.7150 1484.3650 ;
        RECT 99.3850 1487.6350 99.7150 1487.9650 ;
        RECT 99.3850 1491.2350 99.7150 1491.5650 ;
        RECT 99.3850 1494.8350 99.7150 1495.1650 ;
        RECT 99.3850 1498.4350 99.7150 1498.7650 ;
        RECT 99.3850 1502.0350 99.7150 1502.3650 ;
        RECT 99.3850 1505.6350 99.7150 1505.9650 ;
        RECT 99.3850 1509.2350 99.7150 1509.5650 ;
        RECT 99.3850 1512.8350 99.7150 1513.1650 ;
        RECT 99.3850 1516.4350 99.7150 1516.7650 ;
        RECT 99.4100 1520.0350 99.7400 1520.3650 ;
        RECT 920.1200 1012.4350 920.4500 1012.7650 ;
        RECT 920.1200 810.8350 920.4500 811.1650 ;
        RECT 920.1200 814.4350 920.4500 814.7650 ;
        RECT 920.1200 818.0350 920.4500 818.3650 ;
        RECT 920.1200 821.6350 920.4500 821.9650 ;
        RECT 920.1200 828.8350 920.4500 829.1650 ;
        RECT 920.1200 825.2350 920.4500 825.5650 ;
        RECT 920.1200 832.4350 920.4500 832.7650 ;
        RECT 920.1200 836.0350 920.4500 836.3650 ;
        RECT 920.1200 839.6350 920.4500 839.9650 ;
        RECT 920.1200 843.2350 920.4500 843.5650 ;
        RECT 920.1200 846.8350 920.4500 847.1650 ;
        RECT 920.1200 854.0350 920.4500 854.3650 ;
        RECT 920.1200 850.4350 920.4500 850.7650 ;
        RECT 920.1200 857.6350 920.4500 857.9650 ;
        RECT 920.1200 861.2350 920.4500 861.5650 ;
        RECT 920.1200 864.8350 920.4500 865.1650 ;
        RECT 920.1200 868.4350 920.4500 868.7650 ;
        RECT 920.1200 872.0350 920.4500 872.3650 ;
        RECT 920.1200 875.6350 920.4500 875.9650 ;
        RECT 920.1200 879.2350 920.4500 879.5650 ;
        RECT 920.1200 882.8350 920.4500 883.1650 ;
        RECT 920.1200 886.4350 920.4500 886.7650 ;
        RECT 920.1200 890.0350 920.4500 890.3650 ;
        RECT 920.1200 893.6350 920.4500 893.9650 ;
        RECT 920.1200 897.2350 920.4500 897.5650 ;
        RECT 920.1200 900.8350 920.4500 901.1650 ;
        RECT 920.1200 904.4350 920.4500 904.7650 ;
        RECT 920.1200 908.0350 920.4500 908.3650 ;
        RECT 920.1200 911.6350 920.4500 911.9650 ;
        RECT 920.1200 915.2350 920.4500 915.5650 ;
        RECT 920.1200 918.8350 920.4500 919.1650 ;
        RECT 920.1200 922.4350 920.4500 922.7650 ;
        RECT 920.1200 926.0350 920.4500 926.3650 ;
        RECT 920.1200 929.6350 920.4500 929.9650 ;
        RECT 920.1200 933.2350 920.4500 933.5650 ;
        RECT 920.1200 936.8350 920.4500 937.1650 ;
        RECT 920.1200 940.4350 920.4500 940.7650 ;
        RECT 920.1200 944.0350 920.4500 944.3650 ;
        RECT 920.1200 947.6350 920.4500 947.9650 ;
        RECT 920.1200 951.2350 920.4500 951.5650 ;
        RECT 920.1200 954.8350 920.4500 955.1650 ;
        RECT 920.1200 958.4350 920.4500 958.7650 ;
        RECT 920.1200 962.0350 920.4500 962.3650 ;
        RECT 920.1200 965.6350 920.4500 965.9650 ;
        RECT 920.1200 969.2350 920.4500 969.5650 ;
        RECT 920.1200 972.8350 920.4500 973.1650 ;
        RECT 920.1200 976.4350 920.4500 976.7650 ;
        RECT 920.1200 980.0350 920.4500 980.3650 ;
        RECT 920.1200 983.6350 920.4500 983.9650 ;
        RECT 920.1200 987.2350 920.4500 987.5650 ;
        RECT 920.1200 990.8350 920.4500 991.1650 ;
        RECT 920.1200 994.4350 920.4500 994.7650 ;
        RECT 920.1200 998.0350 920.4500 998.3650 ;
        RECT 920.1200 1005.2350 920.4500 1005.5650 ;
        RECT 920.1200 1001.6350 920.4500 1001.9650 ;
        RECT 920.1200 1008.8350 920.4500 1009.1650 ;
        RECT 920.1200 1016.0350 920.4500 1016.3650 ;
        RECT 920.1200 1019.6350 920.4500 1019.9650 ;
        RECT 920.1200 1102.4350 920.4500 1102.7650 ;
        RECT 920.1200 1106.0350 920.4500 1106.3650 ;
        RECT 920.1200 1109.6350 920.4500 1109.9650 ;
        RECT 920.1200 1113.2350 920.4500 1113.5650 ;
        RECT 920.1200 1116.8350 920.4500 1117.1650 ;
        RECT 920.1200 1120.4350 920.4500 1120.7650 ;
        RECT 920.1200 1124.0350 920.4500 1124.3650 ;
        RECT 920.1200 1127.6350 920.4500 1127.9650 ;
        RECT 920.1200 1131.2350 920.4500 1131.5650 ;
        RECT 920.1200 1134.8350 920.4500 1135.1650 ;
        RECT 920.1200 1138.4350 920.4500 1138.7650 ;
        RECT 920.1200 1142.0350 920.4500 1142.3650 ;
        RECT 920.1200 1145.6350 920.4500 1145.9650 ;
        RECT 920.1200 1149.2350 920.4500 1149.5650 ;
        RECT 920.1200 1152.8350 920.4500 1153.1650 ;
        RECT 920.1200 1156.4350 920.4500 1156.7650 ;
        RECT 920.1200 1160.0350 920.4500 1160.3650 ;
        RECT 920.1200 1163.6350 920.4500 1163.9650 ;
        RECT 920.1200 1167.2350 920.4500 1167.5650 ;
        RECT 920.1200 1170.8350 920.4500 1171.1650 ;
        RECT 920.1200 1174.4350 920.4500 1174.7650 ;
        RECT 920.1200 1178.0350 920.4500 1178.3650 ;
        RECT 920.1200 1181.6350 920.4500 1181.9650 ;
        RECT 920.1200 1185.2350 920.4500 1185.5650 ;
        RECT 920.1200 1188.8350 920.4500 1189.1650 ;
        RECT 920.1200 1192.4350 920.4500 1192.7650 ;
        RECT 920.1200 1196.0350 920.4500 1196.3650 ;
        RECT 920.1200 1199.6350 920.4500 1199.9650 ;
        RECT 920.1200 1203.2350 920.4500 1203.5650 ;
        RECT 920.1200 1206.8350 920.4500 1207.1650 ;
        RECT 920.1200 1210.4350 920.4500 1210.7650 ;
        RECT 920.1200 1214.0350 920.4500 1214.3650 ;
        RECT 920.1200 1221.2350 920.4500 1221.5650 ;
        RECT 920.1200 1217.6350 920.4500 1217.9650 ;
        RECT 920.1200 1224.8350 920.4500 1225.1650 ;
        RECT 920.1200 1228.4350 920.4500 1228.7650 ;
        RECT 920.1200 1232.0350 920.4500 1232.3650 ;
        RECT 920.1200 1235.6350 920.4500 1235.9650 ;
        RECT 920.1200 1239.2350 920.4500 1239.5650 ;
        RECT 920.1200 1246.4350 920.4500 1246.7650 ;
        RECT 920.1200 1242.8350 920.4500 1243.1650 ;
        RECT 920.1200 1250.0350 920.4500 1250.3650 ;
        RECT 920.1200 1253.6350 920.4500 1253.9650 ;
        RECT 920.1200 1257.2350 920.4500 1257.5650 ;
        RECT 920.1200 1260.8350 920.4500 1261.1650 ;
        RECT 920.1200 1264.4350 920.4500 1264.7650 ;
        RECT 920.1200 1271.6350 920.4500 1271.9650 ;
        RECT 920.1200 1268.0350 920.4500 1268.3650 ;
        RECT 920.1200 1275.2350 920.4500 1275.5650 ;
        RECT 920.1200 1278.8350 920.4500 1279.1650 ;
        RECT 920.1200 1282.4350 920.4500 1282.7650 ;
        RECT 920.1200 1286.0350 920.4500 1286.3650 ;
        RECT 920.1200 1289.6350 920.4500 1289.9650 ;
        RECT 920.1200 1293.2350 920.4500 1293.5650 ;
        RECT 920.1200 1296.8350 920.4500 1297.1650 ;
        RECT 920.1200 1300.4350 920.4500 1300.7650 ;
        RECT 920.1200 1304.0350 920.4500 1304.3650 ;
        RECT 920.1200 1307.6350 920.4500 1307.9650 ;
        RECT 920.1200 1311.2350 920.4500 1311.5650 ;
        RECT 920.1200 1314.8350 920.4500 1315.1650 ;
        RECT 920.1200 1318.4350 920.4500 1318.7650 ;
        RECT 920.1200 1322.0350 920.4500 1322.3650 ;
        RECT 920.1200 1325.6350 920.4500 1325.9650 ;
        RECT 920.1200 1329.2350 920.4500 1329.5650 ;
        RECT 920.1200 1332.8350 920.4500 1333.1650 ;
        RECT 920.1200 1336.4350 920.4500 1336.7650 ;
        RECT 920.1200 1340.0350 920.4500 1340.3650 ;
        RECT 920.1200 1343.6350 920.4500 1343.9650 ;
        RECT 920.1200 1347.2350 920.4500 1347.5650 ;
        RECT 920.1200 1350.8350 920.4500 1351.1650 ;
        RECT 920.1200 1354.4350 920.4500 1354.7650 ;
        RECT 920.1200 1358.0350 920.4500 1358.3650 ;
        RECT 920.1200 1361.6350 920.4500 1361.9650 ;
        RECT 920.1200 1365.2350 920.4500 1365.5650 ;
        RECT 920.1200 1368.8350 920.4500 1369.1650 ;
        RECT 920.1200 1372.4350 920.4500 1372.7650 ;
        RECT 920.1200 1376.0350 920.4500 1376.3650 ;
        RECT 920.1200 1379.6350 920.4500 1379.9650 ;
        RECT 920.1200 1383.2350 920.4500 1383.5650 ;
        RECT 920.1200 1386.8350 920.4500 1387.1650 ;
        RECT 920.1200 1390.4350 920.4500 1390.7650 ;
        RECT 920.1200 1404.8350 920.4500 1405.1650 ;
        RECT 920.1200 1394.0350 920.4500 1394.3650 ;
        RECT 920.1200 1397.6350 920.4500 1397.9650 ;
        RECT 920.1200 1401.2350 920.4500 1401.5650 ;
        RECT 920.1200 1408.4350 920.4500 1408.7650 ;
        RECT 920.1200 1412.0350 920.4500 1412.3650 ;
        RECT 920.1200 1415.6350 920.4500 1415.9650 ;
        RECT 920.1200 1430.0350 920.4500 1430.3650 ;
        RECT 920.1200 1422.8350 920.4500 1423.1650 ;
        RECT 920.1200 1419.2350 920.4500 1419.5650 ;
        RECT 920.1200 1426.4350 920.4500 1426.7650 ;
        RECT 920.1200 1433.6350 920.4500 1433.9650 ;
        RECT 920.1200 1437.2350 920.4500 1437.5650 ;
        RECT 920.1200 1440.8350 920.4500 1441.1650 ;
        RECT 920.1200 1455.2350 920.4500 1455.5650 ;
        RECT 920.1200 1448.0350 920.4500 1448.3650 ;
        RECT 920.1200 1444.4350 920.4500 1444.7650 ;
        RECT 920.1200 1451.6350 920.4500 1451.9650 ;
        RECT 920.1200 1458.8350 920.4500 1459.1650 ;
        RECT 920.1200 1462.4350 920.4500 1462.7650 ;
        RECT 920.1200 1466.0350 920.4500 1466.3650 ;
        RECT 920.1200 1469.6350 920.4500 1469.9650 ;
        RECT 920.1200 1473.2350 920.4500 1473.5650 ;
        RECT 920.1200 1476.8350 920.4500 1477.1650 ;
        RECT 920.1200 1480.4350 920.4500 1480.7650 ;
        RECT 920.1200 1484.0350 920.4500 1484.3650 ;
        RECT 920.1200 1487.6350 920.4500 1487.9650 ;
        RECT 920.1200 1491.2350 920.4500 1491.5650 ;
        RECT 920.1200 1494.8350 920.4500 1495.1650 ;
        RECT 920.1200 1498.4350 920.4500 1498.7650 ;
        RECT 920.1200 1502.0350 920.4500 1502.3650 ;
        RECT 920.1200 1505.6350 920.4500 1505.9650 ;
        RECT 920.1200 1509.2350 920.4500 1509.5650 ;
        RECT 920.1200 1512.8350 920.4500 1513.1650 ;
        RECT 920.1200 1516.4350 920.4500 1516.7650 ;
        RECT 920.0950 1520.0350 920.4250 1520.3650 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 110.0000 610.0000 111.0000 1010.0000 ;
        RECT 223.8550 610.0000 224.8550 1010.0000 ;
        RECT 337.7100 610.0000 338.7100 1010.0000 ;
        RECT 451.5650 610.0000 452.5650 1010.0000 ;
        RECT 565.4200 610.0000 566.4200 1010.0000 ;
        RECT 679.2750 610.0000 680.2750 1010.0000 ;
        RECT 793.1300 610.0000 794.1300 1010.0000 ;
        RECT 906.9850 610.0000 907.9850 1010.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 110.0000 1110.0000 111.0000 1510.0000 ;
        RECT 223.8550 1110.0000 224.8550 1510.0000 ;
        RECT 337.7100 1110.0000 338.7100 1510.0000 ;
        RECT 451.5650 1110.0000 452.5650 1510.0000 ;
        RECT 565.4200 1110.0000 566.4200 1510.0000 ;
        RECT 679.2750 1110.0000 680.2750 1510.0000 ;
        RECT 793.1300 1110.0000 794.1300 1510.0000 ;
        RECT 906.9850 1110.0000 907.9850 1510.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 110.0000 110.0000 111.0000 510.0000 ;
        RECT 223.8550 110.0000 224.8550 510.0000 ;
        RECT 337.7100 110.0000 338.7100 510.0000 ;
        RECT 451.5650 110.0000 452.5650 510.0000 ;
        RECT 565.4200 110.0000 566.4200 510.0000 ;
        RECT 679.2750 110.0000 680.2750 510.0000 ;
        RECT 793.1300 110.0000 794.1300 510.0000 ;
        RECT 906.9850 110.0000 907.9850 510.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 1008.0000 10.0000 1010.0000 1610.0000 ;
        RECT 898.0000 10.0000 900.0000 1610.0000 ;
        RECT 788.0000 10.0000 790.0000 1610.0000 ;
        RECT 678.0000 10.0000 680.0000 1610.0000 ;
        RECT 568.0000 10.0000 570.0000 1610.0000 ;
        RECT 458.0000 10.0000 460.0000 1610.0000 ;
        RECT 348.0000 10.0000 350.0000 1610.0000 ;
        RECT 238.0000 10.0000 240.0000 1610.0000 ;
        RECT 128.0000 10.0000 130.0000 1610.0000 ;
        RECT 18.0000 10.0000 20.0000 1610.0000 ;
        RECT 18.0000 9.8350 20.0000 10.1650 ;
        RECT 128.0000 9.8350 130.0000 10.1650 ;
        RECT 238.0000 9.8350 240.0000 10.1650 ;
        RECT 348.0000 9.8350 350.0000 10.1650 ;
        RECT 458.0000 9.8350 460.0000 10.1650 ;
        RECT 568.0000 9.8350 570.0000 10.1650 ;
        RECT 678.0000 9.8350 680.0000 10.1650 ;
        RECT 788.0000 9.8350 790.0000 10.1650 ;
        RECT 898.0000 9.8350 900.0000 10.1650 ;
        RECT 1008.0000 9.8350 1010.0000 10.1650 ;
        RECT 99.3850 99.8350 99.7150 100.1650 ;
        RECT 99.3850 103.4350 99.7150 103.7650 ;
        RECT 99.3850 107.0350 99.7150 107.3650 ;
        RECT 99.3850 110.6350 99.7150 110.9650 ;
        RECT 99.3850 114.2350 99.7150 114.5650 ;
        RECT 99.3850 117.8350 99.7150 118.1650 ;
        RECT 99.3850 121.4350 99.7150 121.7650 ;
        RECT 99.3850 125.0350 99.7150 125.3650 ;
        RECT 99.3850 128.6350 99.7150 128.9650 ;
        RECT 99.3850 132.2350 99.7150 132.5650 ;
        RECT 99.3850 135.8350 99.7150 136.1650 ;
        RECT 99.3850 139.4350 99.7150 139.7650 ;
        RECT 99.3850 143.0350 99.7150 143.3650 ;
        RECT 99.3850 146.6350 99.7150 146.9650 ;
        RECT 99.3850 150.2350 99.7150 150.5650 ;
        RECT 99.3850 153.8350 99.7150 154.1650 ;
        RECT 99.3850 157.4350 99.7150 157.7650 ;
        RECT 99.3850 161.0350 99.7150 161.3650 ;
        RECT 99.3850 164.6350 99.7150 164.9650 ;
        RECT 99.3850 168.2350 99.7150 168.5650 ;
        RECT 99.3850 171.8350 99.7150 172.1650 ;
        RECT 99.3850 175.4350 99.7150 175.7650 ;
        RECT 99.3850 189.8350 99.7150 190.1650 ;
        RECT 99.3850 179.0350 99.7150 179.3650 ;
        RECT 99.3850 182.6350 99.7150 182.9650 ;
        RECT 99.3850 186.2350 99.7150 186.5650 ;
        RECT 99.3850 193.4350 99.7150 193.7650 ;
        RECT 99.3850 197.0350 99.7150 197.3650 ;
        RECT 99.3850 200.6350 99.7150 200.9650 ;
        RECT 99.3850 215.0350 99.7150 215.3650 ;
        RECT 99.3850 204.2350 99.7150 204.5650 ;
        RECT 99.3850 207.8350 99.7150 208.1650 ;
        RECT 99.3850 211.4350 99.7150 211.7650 ;
        RECT 99.3850 218.6350 99.7150 218.9650 ;
        RECT 99.3850 222.2350 99.7150 222.5650 ;
        RECT 99.3850 225.8350 99.7150 226.1650 ;
        RECT 99.3850 240.2350 99.7150 240.5650 ;
        RECT 99.3850 229.4350 99.7150 229.7650 ;
        RECT 99.3850 233.0350 99.7150 233.3650 ;
        RECT 99.3850 236.6350 99.7150 236.9650 ;
        RECT 99.3850 243.8350 99.7150 244.1650 ;
        RECT 99.3850 247.4350 99.7150 247.7650 ;
        RECT 99.3850 251.0350 99.7150 251.3650 ;
        RECT 99.3850 254.6350 99.7150 254.9650 ;
        RECT 99.3850 258.2350 99.7150 258.5650 ;
        RECT 99.3850 261.8350 99.7150 262.1650 ;
        RECT 99.3850 265.4350 99.7150 265.7650 ;
        RECT 99.3850 269.0350 99.7150 269.3650 ;
        RECT 99.3850 272.6350 99.7150 272.9650 ;
        RECT 99.3850 276.2350 99.7150 276.5650 ;
        RECT 99.3850 279.8350 99.7150 280.1650 ;
        RECT 99.3850 283.4350 99.7150 283.7650 ;
        RECT 99.3850 287.0350 99.7150 287.3650 ;
        RECT 99.3850 290.6350 99.7150 290.9650 ;
        RECT 99.3850 294.2350 99.7150 294.5650 ;
        RECT 99.3850 297.8350 99.7150 298.1650 ;
        RECT 99.3850 301.4350 99.7150 301.7650 ;
        RECT 99.3850 305.0350 99.7150 305.3650 ;
        RECT 99.3850 308.6350 99.7150 308.9650 ;
        RECT 99.3850 312.2350 99.7150 312.5650 ;
        RECT 99.3850 315.8350 99.7150 316.1650 ;
        RECT 99.3850 319.4350 99.7150 319.7650 ;
        RECT 99.3850 323.0350 99.7150 323.3650 ;
        RECT 99.3850 326.6350 99.7150 326.9650 ;
        RECT 99.3850 330.2350 99.7150 330.5650 ;
        RECT 99.3850 333.8350 99.7150 334.1650 ;
        RECT 99.3850 337.4350 99.7150 337.7650 ;
        RECT 99.3850 341.0350 99.7150 341.3650 ;
        RECT 99.3850 344.6350 99.7150 344.9650 ;
        RECT 99.3850 348.2350 99.7150 348.5650 ;
        RECT 99.3850 351.8350 99.7150 352.1650 ;
        RECT 99.3850 355.4350 99.7150 355.7650 ;
        RECT 99.3850 359.0350 99.7150 359.3650 ;
        RECT 99.3850 362.6350 99.7150 362.9650 ;
        RECT 99.3850 366.2350 99.7150 366.5650 ;
        RECT 99.3850 369.8350 99.7150 370.1650 ;
        RECT 99.3850 373.4350 99.7150 373.7650 ;
        RECT 99.3850 377.0350 99.7150 377.3650 ;
        RECT 99.3850 380.6350 99.7150 380.9650 ;
        RECT 99.3850 384.2350 99.7150 384.5650 ;
        RECT 99.3850 387.8350 99.7150 388.1650 ;
        RECT 99.3850 391.4350 99.7150 391.7650 ;
        RECT 99.3850 398.6350 99.7150 398.9650 ;
        RECT 99.3850 395.0350 99.7150 395.3650 ;
        RECT 99.3850 402.2350 99.7150 402.5650 ;
        RECT 99.3850 607.4350 99.7150 607.7650 ;
        RECT 99.3850 405.8350 99.7150 406.1650 ;
        RECT 99.3850 409.4350 99.7150 409.7650 ;
        RECT 99.3850 413.0350 99.7150 413.3650 ;
        RECT 99.3850 416.6350 99.7150 416.9650 ;
        RECT 99.3850 423.8350 99.7150 424.1650 ;
        RECT 99.3850 420.2350 99.7150 420.5650 ;
        RECT 99.3850 427.4350 99.7150 427.7650 ;
        RECT 99.3850 431.0350 99.7150 431.3650 ;
        RECT 99.3850 434.6350 99.7150 434.9650 ;
        RECT 99.3850 438.2350 99.7150 438.5650 ;
        RECT 99.3850 441.8350 99.7150 442.1650 ;
        RECT 99.3850 449.0350 99.7150 449.3650 ;
        RECT 99.3850 445.4350 99.7150 445.7650 ;
        RECT 99.3850 452.6350 99.7150 452.9650 ;
        RECT 99.3850 456.2350 99.7150 456.5650 ;
        RECT 99.3850 459.8350 99.7150 460.1650 ;
        RECT 99.3850 463.4350 99.7150 463.7650 ;
        RECT 99.3850 467.0350 99.7150 467.3650 ;
        RECT 99.3850 470.6350 99.7150 470.9650 ;
        RECT 99.3850 474.2350 99.7150 474.5650 ;
        RECT 99.3850 477.8350 99.7150 478.1650 ;
        RECT 99.3850 481.4350 99.7150 481.7650 ;
        RECT 99.3850 485.0350 99.7150 485.3650 ;
        RECT 99.3850 488.6350 99.7150 488.9650 ;
        RECT 99.3850 492.2350 99.7150 492.5650 ;
        RECT 99.3850 495.8350 99.7150 496.1650 ;
        RECT 99.3850 499.4350 99.7150 499.7650 ;
        RECT 99.3850 503.0350 99.7150 503.3650 ;
        RECT 99.3850 506.6350 99.7150 506.9650 ;
        RECT 99.3850 510.2350 99.7150 510.5650 ;
        RECT 99.3850 513.8350 99.7150 514.1650 ;
        RECT 99.3850 517.4350 99.7150 517.7650 ;
        RECT 99.3850 600.2350 99.7150 600.5650 ;
        RECT 99.3850 603.8350 99.7150 604.1650 ;
        RECT 99.3850 657.8350 99.7150 658.1650 ;
        RECT 99.3850 632.6350 99.7150 632.9650 ;
        RECT 99.3850 611.0350 99.7150 611.3650 ;
        RECT 99.3850 614.6350 99.7150 614.9650 ;
        RECT 99.3850 618.2350 99.7150 618.5650 ;
        RECT 99.3850 621.8350 99.7150 622.1650 ;
        RECT 99.3850 625.4350 99.7150 625.7650 ;
        RECT 99.3850 629.0350 99.7150 629.3650 ;
        RECT 99.3850 636.2350 99.7150 636.5650 ;
        RECT 99.3850 639.8350 99.7150 640.1650 ;
        RECT 99.3850 643.4350 99.7150 643.7650 ;
        RECT 99.3850 647.0350 99.7150 647.3650 ;
        RECT 99.3850 650.6350 99.7150 650.9650 ;
        RECT 99.3850 654.2350 99.7150 654.5650 ;
        RECT 99.3850 661.4350 99.7150 661.7650 ;
        RECT 99.3850 665.0350 99.7150 665.3650 ;
        RECT 99.3850 668.6350 99.7150 668.9650 ;
        RECT 99.3850 672.2350 99.7150 672.5650 ;
        RECT 99.3850 675.8350 99.7150 676.1650 ;
        RECT 99.3850 679.4350 99.7150 679.7650 ;
        RECT 99.3850 683.0350 99.7150 683.3650 ;
        RECT 99.3850 686.6350 99.7150 686.9650 ;
        RECT 99.3850 690.2350 99.7150 690.5650 ;
        RECT 99.3850 693.8350 99.7150 694.1650 ;
        RECT 99.3850 697.4350 99.7150 697.7650 ;
        RECT 99.3850 701.0350 99.7150 701.3650 ;
        RECT 99.3850 704.6350 99.7150 704.9650 ;
        RECT 99.3850 708.2350 99.7150 708.5650 ;
        RECT 99.3850 711.8350 99.7150 712.1650 ;
        RECT 99.3850 715.4350 99.7150 715.7650 ;
        RECT 99.3850 719.0350 99.7150 719.3650 ;
        RECT 99.3850 722.6350 99.7150 722.9650 ;
        RECT 99.3850 726.2350 99.7150 726.5650 ;
        RECT 99.3850 729.8350 99.7150 730.1650 ;
        RECT 99.3850 733.4350 99.7150 733.7650 ;
        RECT 99.3850 737.0350 99.7150 737.3650 ;
        RECT 99.3850 740.6350 99.7150 740.9650 ;
        RECT 99.3850 744.2350 99.7150 744.5650 ;
        RECT 99.3850 747.8350 99.7150 748.1650 ;
        RECT 99.3850 751.4350 99.7150 751.7650 ;
        RECT 99.3850 755.0350 99.7150 755.3650 ;
        RECT 99.3850 758.6350 99.7150 758.9650 ;
        RECT 99.3850 762.2350 99.7150 762.5650 ;
        RECT 99.3850 765.8350 99.7150 766.1650 ;
        RECT 99.3850 769.4350 99.7150 769.7650 ;
        RECT 99.3850 773.0350 99.7150 773.3650 ;
        RECT 99.3850 776.6350 99.7150 776.9650 ;
        RECT 99.3850 780.2350 99.7150 780.5650 ;
        RECT 99.3850 783.8350 99.7150 784.1650 ;
        RECT 99.3850 787.4350 99.7150 787.7650 ;
        RECT 99.3850 791.0350 99.7150 791.3650 ;
        RECT 99.3850 794.6350 99.7150 794.9650 ;
        RECT 99.3850 798.2350 99.7150 798.5650 ;
        RECT 99.3850 801.8350 99.7150 802.1650 ;
        RECT 99.3850 805.4350 99.7150 805.7650 ;
        RECT 99.3850 809.0350 99.7150 809.3650 ;
        RECT 920.1200 99.8350 920.4500 100.1650 ;
        RECT 920.1200 103.4350 920.4500 103.7650 ;
        RECT 920.1200 107.0350 920.4500 107.3650 ;
        RECT 920.1200 110.6350 920.4500 110.9650 ;
        RECT 920.1200 114.2350 920.4500 114.5650 ;
        RECT 920.1200 117.8350 920.4500 118.1650 ;
        RECT 920.1200 121.4350 920.4500 121.7650 ;
        RECT 920.1200 125.0350 920.4500 125.3650 ;
        RECT 920.1200 128.6350 920.4500 128.9650 ;
        RECT 920.1200 132.2350 920.4500 132.5650 ;
        RECT 920.1200 135.8350 920.4500 136.1650 ;
        RECT 920.1200 139.4350 920.4500 139.7650 ;
        RECT 920.1200 143.0350 920.4500 143.3650 ;
        RECT 920.1200 146.6350 920.4500 146.9650 ;
        RECT 920.1200 150.2350 920.4500 150.5650 ;
        RECT 920.1200 153.8350 920.4500 154.1650 ;
        RECT 920.1200 157.4350 920.4500 157.7650 ;
        RECT 920.1200 161.0350 920.4500 161.3650 ;
        RECT 920.1200 164.6350 920.4500 164.9650 ;
        RECT 920.1200 168.2350 920.4500 168.5650 ;
        RECT 920.1200 171.8350 920.4500 172.1650 ;
        RECT 920.1200 175.4350 920.4500 175.7650 ;
        RECT 920.1200 189.8350 920.4500 190.1650 ;
        RECT 920.1200 179.0350 920.4500 179.3650 ;
        RECT 920.1200 182.6350 920.4500 182.9650 ;
        RECT 920.1200 186.2350 920.4500 186.5650 ;
        RECT 920.1200 193.4350 920.4500 193.7650 ;
        RECT 920.1200 197.0350 920.4500 197.3650 ;
        RECT 920.1200 200.6350 920.4500 200.9650 ;
        RECT 920.1200 215.0350 920.4500 215.3650 ;
        RECT 920.1200 204.2350 920.4500 204.5650 ;
        RECT 920.1200 207.8350 920.4500 208.1650 ;
        RECT 920.1200 211.4350 920.4500 211.7650 ;
        RECT 920.1200 218.6350 920.4500 218.9650 ;
        RECT 920.1200 222.2350 920.4500 222.5650 ;
        RECT 920.1200 225.8350 920.4500 226.1650 ;
        RECT 920.1200 240.2350 920.4500 240.5650 ;
        RECT 920.1200 229.4350 920.4500 229.7650 ;
        RECT 920.1200 233.0350 920.4500 233.3650 ;
        RECT 920.1200 236.6350 920.4500 236.9650 ;
        RECT 920.1200 243.8350 920.4500 244.1650 ;
        RECT 920.1200 247.4350 920.4500 247.7650 ;
        RECT 920.1200 251.0350 920.4500 251.3650 ;
        RECT 920.1200 254.6350 920.4500 254.9650 ;
        RECT 920.1200 258.2350 920.4500 258.5650 ;
        RECT 920.1200 261.8350 920.4500 262.1650 ;
        RECT 920.1200 265.4350 920.4500 265.7650 ;
        RECT 920.1200 269.0350 920.4500 269.3650 ;
        RECT 920.1200 272.6350 920.4500 272.9650 ;
        RECT 920.1200 276.2350 920.4500 276.5650 ;
        RECT 920.1200 279.8350 920.4500 280.1650 ;
        RECT 920.1200 283.4350 920.4500 283.7650 ;
        RECT 920.1200 287.0350 920.4500 287.3650 ;
        RECT 920.1200 290.6350 920.4500 290.9650 ;
        RECT 920.1200 294.2350 920.4500 294.5650 ;
        RECT 920.1200 297.8350 920.4500 298.1650 ;
        RECT 920.1200 301.4350 920.4500 301.7650 ;
        RECT 920.1200 305.0350 920.4500 305.3650 ;
        RECT 920.1200 308.6350 920.4500 308.9650 ;
        RECT 920.1200 312.2350 920.4500 312.5650 ;
        RECT 920.1200 315.8350 920.4500 316.1650 ;
        RECT 920.1200 319.4350 920.4500 319.7650 ;
        RECT 920.1200 323.0350 920.4500 323.3650 ;
        RECT 920.1200 326.6350 920.4500 326.9650 ;
        RECT 920.1200 330.2350 920.4500 330.5650 ;
        RECT 920.1200 333.8350 920.4500 334.1650 ;
        RECT 920.1200 337.4350 920.4500 337.7650 ;
        RECT 920.1200 341.0350 920.4500 341.3650 ;
        RECT 920.1200 344.6350 920.4500 344.9650 ;
        RECT 920.1200 348.2350 920.4500 348.5650 ;
        RECT 920.1200 351.8350 920.4500 352.1650 ;
        RECT 920.1200 355.4350 920.4500 355.7650 ;
        RECT 920.1200 359.0350 920.4500 359.3650 ;
        RECT 920.1200 362.6350 920.4500 362.9650 ;
        RECT 920.1200 366.2350 920.4500 366.5650 ;
        RECT 920.1200 369.8350 920.4500 370.1650 ;
        RECT 920.1200 373.4350 920.4500 373.7650 ;
        RECT 920.1200 377.0350 920.4500 377.3650 ;
        RECT 920.1200 380.6350 920.4500 380.9650 ;
        RECT 920.1200 384.2350 920.4500 384.5650 ;
        RECT 920.1200 387.8350 920.4500 388.1650 ;
        RECT 920.1200 391.4350 920.4500 391.7650 ;
        RECT 920.1200 398.6350 920.4500 398.9650 ;
        RECT 920.1200 395.0350 920.4500 395.3650 ;
        RECT 920.1200 402.2350 920.4500 402.5650 ;
        RECT 920.1200 607.4350 920.4500 607.7650 ;
        RECT 920.1200 405.8350 920.4500 406.1650 ;
        RECT 920.1200 409.4350 920.4500 409.7650 ;
        RECT 920.1200 413.0350 920.4500 413.3650 ;
        RECT 920.1200 416.6350 920.4500 416.9650 ;
        RECT 920.1200 423.8350 920.4500 424.1650 ;
        RECT 920.1200 420.2350 920.4500 420.5650 ;
        RECT 920.1200 427.4350 920.4500 427.7650 ;
        RECT 920.1200 431.0350 920.4500 431.3650 ;
        RECT 920.1200 434.6350 920.4500 434.9650 ;
        RECT 920.1200 438.2350 920.4500 438.5650 ;
        RECT 920.1200 441.8350 920.4500 442.1650 ;
        RECT 920.1200 449.0350 920.4500 449.3650 ;
        RECT 920.1200 445.4350 920.4500 445.7650 ;
        RECT 920.1200 452.6350 920.4500 452.9650 ;
        RECT 920.1200 456.2350 920.4500 456.5650 ;
        RECT 920.1200 459.8350 920.4500 460.1650 ;
        RECT 920.1200 463.4350 920.4500 463.7650 ;
        RECT 920.1200 467.0350 920.4500 467.3650 ;
        RECT 920.1200 470.6350 920.4500 470.9650 ;
        RECT 920.1200 474.2350 920.4500 474.5650 ;
        RECT 920.1200 477.8350 920.4500 478.1650 ;
        RECT 920.1200 481.4350 920.4500 481.7650 ;
        RECT 920.1200 485.0350 920.4500 485.3650 ;
        RECT 920.1200 488.6350 920.4500 488.9650 ;
        RECT 920.1200 492.2350 920.4500 492.5650 ;
        RECT 920.1200 495.8350 920.4500 496.1650 ;
        RECT 920.1200 499.4350 920.4500 499.7650 ;
        RECT 920.1200 503.0350 920.4500 503.3650 ;
        RECT 920.1200 506.6350 920.4500 506.9650 ;
        RECT 920.1200 510.2350 920.4500 510.5650 ;
        RECT 920.1200 513.8350 920.4500 514.1650 ;
        RECT 920.1200 517.4350 920.4500 517.7650 ;
        RECT 920.1200 600.2350 920.4500 600.5650 ;
        RECT 920.1200 603.8350 920.4500 604.1650 ;
        RECT 920.1200 657.8350 920.4500 658.1650 ;
        RECT 920.1200 632.6350 920.4500 632.9650 ;
        RECT 920.1200 611.0350 920.4500 611.3650 ;
        RECT 920.1200 614.6350 920.4500 614.9650 ;
        RECT 920.1200 618.2350 920.4500 618.5650 ;
        RECT 920.1200 621.8350 920.4500 622.1650 ;
        RECT 920.1200 625.4350 920.4500 625.7650 ;
        RECT 920.1200 629.0350 920.4500 629.3650 ;
        RECT 920.1200 636.2350 920.4500 636.5650 ;
        RECT 920.1200 639.8350 920.4500 640.1650 ;
        RECT 920.1200 643.4350 920.4500 643.7650 ;
        RECT 920.1200 647.0350 920.4500 647.3650 ;
        RECT 920.1200 650.6350 920.4500 650.9650 ;
        RECT 920.1200 654.2350 920.4500 654.5650 ;
        RECT 920.1200 661.4350 920.4500 661.7650 ;
        RECT 920.1200 665.0350 920.4500 665.3650 ;
        RECT 920.1200 668.6350 920.4500 668.9650 ;
        RECT 920.1200 672.2350 920.4500 672.5650 ;
        RECT 920.1200 675.8350 920.4500 676.1650 ;
        RECT 920.1200 679.4350 920.4500 679.7650 ;
        RECT 920.1200 683.0350 920.4500 683.3650 ;
        RECT 920.1200 686.6350 920.4500 686.9650 ;
        RECT 920.1200 690.2350 920.4500 690.5650 ;
        RECT 920.1200 693.8350 920.4500 694.1650 ;
        RECT 920.1200 697.4350 920.4500 697.7650 ;
        RECT 920.1200 701.0350 920.4500 701.3650 ;
        RECT 920.1200 704.6350 920.4500 704.9650 ;
        RECT 920.1200 708.2350 920.4500 708.5650 ;
        RECT 920.1200 711.8350 920.4500 712.1650 ;
        RECT 920.1200 715.4350 920.4500 715.7650 ;
        RECT 920.1200 719.0350 920.4500 719.3650 ;
        RECT 920.1200 722.6350 920.4500 722.9650 ;
        RECT 920.1200 726.2350 920.4500 726.5650 ;
        RECT 920.1200 729.8350 920.4500 730.1650 ;
        RECT 920.1200 733.4350 920.4500 733.7650 ;
        RECT 920.1200 737.0350 920.4500 737.3650 ;
        RECT 920.1200 740.6350 920.4500 740.9650 ;
        RECT 920.1200 744.2350 920.4500 744.5650 ;
        RECT 920.1200 747.8350 920.4500 748.1650 ;
        RECT 920.1200 751.4350 920.4500 751.7650 ;
        RECT 920.1200 755.0350 920.4500 755.3650 ;
        RECT 920.1200 758.6350 920.4500 758.9650 ;
        RECT 920.1200 762.2350 920.4500 762.5650 ;
        RECT 920.1200 765.8350 920.4500 766.1650 ;
        RECT 920.1200 769.4350 920.4500 769.7650 ;
        RECT 920.1200 773.0350 920.4500 773.3650 ;
        RECT 920.1200 776.6350 920.4500 776.9650 ;
        RECT 920.1200 780.2350 920.4500 780.5650 ;
        RECT 920.1200 783.8350 920.4500 784.1650 ;
        RECT 920.1200 787.4350 920.4500 787.7650 ;
        RECT 920.1200 791.0350 920.4500 791.3650 ;
        RECT 920.1200 794.6350 920.4500 794.9650 ;
        RECT 920.1200 798.2350 920.4500 798.5650 ;
        RECT 920.1200 801.8350 920.4500 802.1650 ;
        RECT 920.1200 805.4350 920.4500 805.7650 ;
        RECT 920.1200 809.0350 920.4500 809.3650 ;
        RECT 99.3850 816.2350 99.7150 816.5650 ;
        RECT 99.3850 812.6350 99.7150 812.9650 ;
        RECT 99.3850 819.8350 99.7150 820.1650 ;
        RECT 99.3850 823.4350 99.7150 823.7650 ;
        RECT 99.3850 827.0350 99.7150 827.3650 ;
        RECT 99.3850 830.6350 99.7150 830.9650 ;
        RECT 99.3850 834.2350 99.7150 834.5650 ;
        RECT 99.3850 841.4350 99.7150 841.7650 ;
        RECT 99.3850 837.8350 99.7150 838.1650 ;
        RECT 99.3850 845.0350 99.7150 845.3650 ;
        RECT 99.3850 848.6350 99.7150 848.9650 ;
        RECT 99.3850 852.2350 99.7150 852.5650 ;
        RECT 99.3850 855.8350 99.7150 856.1650 ;
        RECT 99.3850 859.4350 99.7150 859.7650 ;
        RECT 99.3850 866.6350 99.7150 866.9650 ;
        RECT 99.3850 863.0350 99.7150 863.3650 ;
        RECT 99.3850 870.2350 99.7150 870.5650 ;
        RECT 99.3850 873.8350 99.7150 874.1650 ;
        RECT 99.3850 877.4350 99.7150 877.7650 ;
        RECT 99.3850 881.0350 99.7150 881.3650 ;
        RECT 99.3850 884.6350 99.7150 884.9650 ;
        RECT 99.3850 888.2350 99.7150 888.5650 ;
        RECT 99.3850 891.8350 99.7150 892.1650 ;
        RECT 99.3850 895.4350 99.7150 895.7650 ;
        RECT 99.3850 899.0350 99.7150 899.3650 ;
        RECT 99.3850 902.6350 99.7150 902.9650 ;
        RECT 99.3850 906.2350 99.7150 906.5650 ;
        RECT 99.3850 909.8350 99.7150 910.1650 ;
        RECT 99.3850 913.4350 99.7150 913.7650 ;
        RECT 99.3850 917.0350 99.7150 917.3650 ;
        RECT 99.3850 920.6350 99.7150 920.9650 ;
        RECT 99.3850 924.2350 99.7150 924.5650 ;
        RECT 99.3850 927.8350 99.7150 928.1650 ;
        RECT 99.3850 931.4350 99.7150 931.7650 ;
        RECT 99.3850 935.0350 99.7150 935.3650 ;
        RECT 99.3850 938.6350 99.7150 938.9650 ;
        RECT 99.3850 942.2350 99.7150 942.5650 ;
        RECT 99.3850 945.8350 99.7150 946.1650 ;
        RECT 99.3850 949.4350 99.7150 949.7650 ;
        RECT 99.3850 953.0350 99.7150 953.3650 ;
        RECT 99.3850 956.6350 99.7150 956.9650 ;
        RECT 99.3850 960.2350 99.7150 960.5650 ;
        RECT 99.3850 963.8350 99.7150 964.1650 ;
        RECT 99.3850 967.4350 99.7150 967.7650 ;
        RECT 99.3850 971.0350 99.7150 971.3650 ;
        RECT 99.3850 974.6350 99.7150 974.9650 ;
        RECT 99.3850 978.2350 99.7150 978.5650 ;
        RECT 99.3850 981.8350 99.7150 982.1650 ;
        RECT 99.3850 985.4350 99.7150 985.7650 ;
        RECT 99.3850 999.8350 99.7150 1000.1650 ;
        RECT 99.3850 989.0350 99.7150 989.3650 ;
        RECT 99.3850 992.6350 99.7150 992.9650 ;
        RECT 99.3850 996.2350 99.7150 996.5650 ;
        RECT 99.3850 1003.4350 99.7150 1003.7650 ;
        RECT 99.3850 1007.0350 99.7150 1007.3650 ;
        RECT 99.3850 1010.6350 99.7150 1010.9650 ;
        RECT 99.3850 1014.2350 99.7150 1014.5650 ;
        RECT 99.3850 1017.8350 99.7150 1018.1650 ;
        RECT 99.3850 1100.6350 99.7150 1100.9650 ;
        RECT 99.3850 1104.2350 99.7150 1104.5650 ;
        RECT 99.3850 1107.8350 99.7150 1108.1650 ;
        RECT 99.3850 1111.4350 99.7150 1111.7650 ;
        RECT 99.3850 1115.0350 99.7150 1115.3650 ;
        RECT 99.3850 1118.6350 99.7150 1118.9650 ;
        RECT 99.3850 1122.2350 99.7150 1122.5650 ;
        RECT 99.3850 1125.8350 99.7150 1126.1650 ;
        RECT 99.3850 1129.4350 99.7150 1129.7650 ;
        RECT 99.3850 1133.0350 99.7150 1133.3650 ;
        RECT 99.3850 1136.6350 99.7150 1136.9650 ;
        RECT 99.3850 1140.2350 99.7150 1140.5650 ;
        RECT 99.3850 1143.8350 99.7150 1144.1650 ;
        RECT 99.3850 1147.4350 99.7150 1147.7650 ;
        RECT 99.3850 1151.0350 99.7150 1151.3650 ;
        RECT 99.3850 1154.6350 99.7150 1154.9650 ;
        RECT 99.3850 1158.2350 99.7150 1158.5650 ;
        RECT 99.3850 1161.8350 99.7150 1162.1650 ;
        RECT 99.3850 1165.4350 99.7150 1165.7650 ;
        RECT 99.3850 1169.0350 99.7150 1169.3650 ;
        RECT 99.3850 1172.6350 99.7150 1172.9650 ;
        RECT 99.3850 1176.2350 99.7150 1176.5650 ;
        RECT 99.3850 1179.8350 99.7150 1180.1650 ;
        RECT 99.3850 1183.4350 99.7150 1183.7650 ;
        RECT 99.3850 1187.0350 99.7150 1187.3650 ;
        RECT 99.3850 1190.6350 99.7150 1190.9650 ;
        RECT 99.3850 1194.2350 99.7150 1194.5650 ;
        RECT 99.3850 1197.8350 99.7150 1198.1650 ;
        RECT 99.3850 1201.4350 99.7150 1201.7650 ;
        RECT 99.3850 1208.6350 99.7150 1208.9650 ;
        RECT 99.3850 1205.0350 99.7150 1205.3650 ;
        RECT 99.3850 1212.2350 99.7150 1212.5650 ;
        RECT 99.3850 1417.4350 99.7150 1417.7650 ;
        RECT 99.3850 1215.8350 99.7150 1216.1650 ;
        RECT 99.3850 1219.4350 99.7150 1219.7650 ;
        RECT 99.3850 1223.0350 99.7150 1223.3650 ;
        RECT 99.3850 1226.6350 99.7150 1226.9650 ;
        RECT 99.3850 1233.8350 99.7150 1234.1650 ;
        RECT 99.3850 1230.2350 99.7150 1230.5650 ;
        RECT 99.3850 1237.4350 99.7150 1237.7650 ;
        RECT 99.3850 1241.0350 99.7150 1241.3650 ;
        RECT 99.3850 1244.6350 99.7150 1244.9650 ;
        RECT 99.3850 1248.2350 99.7150 1248.5650 ;
        RECT 99.3850 1251.8350 99.7150 1252.1650 ;
        RECT 99.3850 1259.0350 99.7150 1259.3650 ;
        RECT 99.3850 1255.4350 99.7150 1255.7650 ;
        RECT 99.3850 1262.6350 99.7150 1262.9650 ;
        RECT 99.3850 1266.2350 99.7150 1266.5650 ;
        RECT 99.3850 1269.8350 99.7150 1270.1650 ;
        RECT 99.3850 1273.4350 99.7150 1273.7650 ;
        RECT 99.3850 1277.0350 99.7150 1277.3650 ;
        RECT 99.3850 1280.6350 99.7150 1280.9650 ;
        RECT 99.3850 1284.2350 99.7150 1284.5650 ;
        RECT 99.3850 1287.8350 99.7150 1288.1650 ;
        RECT 99.3850 1291.4350 99.7150 1291.7650 ;
        RECT 99.3850 1295.0350 99.7150 1295.3650 ;
        RECT 99.3850 1298.6350 99.7150 1298.9650 ;
        RECT 99.3850 1302.2350 99.7150 1302.5650 ;
        RECT 99.3850 1305.8350 99.7150 1306.1650 ;
        RECT 99.3850 1309.4350 99.7150 1309.7650 ;
        RECT 99.3850 1313.0350 99.7150 1313.3650 ;
        RECT 99.3850 1316.6350 99.7150 1316.9650 ;
        RECT 99.3850 1320.2350 99.7150 1320.5650 ;
        RECT 99.3850 1323.8350 99.7150 1324.1650 ;
        RECT 99.3850 1327.4350 99.7150 1327.7650 ;
        RECT 99.3850 1331.0350 99.7150 1331.3650 ;
        RECT 99.3850 1334.6350 99.7150 1334.9650 ;
        RECT 99.3850 1338.2350 99.7150 1338.5650 ;
        RECT 99.3850 1341.8350 99.7150 1342.1650 ;
        RECT 99.3850 1345.4350 99.7150 1345.7650 ;
        RECT 99.3850 1349.0350 99.7150 1349.3650 ;
        RECT 99.3850 1352.6350 99.7150 1352.9650 ;
        RECT 99.3850 1356.2350 99.7150 1356.5650 ;
        RECT 99.3850 1359.8350 99.7150 1360.1650 ;
        RECT 99.3850 1363.4350 99.7150 1363.7650 ;
        RECT 99.3850 1367.0350 99.7150 1367.3650 ;
        RECT 99.3850 1370.6350 99.7150 1370.9650 ;
        RECT 99.3850 1374.2350 99.7150 1374.5650 ;
        RECT 99.3850 1377.8350 99.7150 1378.1650 ;
        RECT 99.3850 1381.4350 99.7150 1381.7650 ;
        RECT 99.3850 1385.0350 99.7150 1385.3650 ;
        RECT 99.3850 1388.6350 99.7150 1388.9650 ;
        RECT 99.3850 1392.2350 99.7150 1392.5650 ;
        RECT 99.3850 1395.8350 99.7150 1396.1650 ;
        RECT 99.3850 1399.4350 99.7150 1399.7650 ;
        RECT 99.3850 1403.0350 99.7150 1403.3650 ;
        RECT 99.3850 1406.6350 99.7150 1406.9650 ;
        RECT 99.3850 1410.2350 99.7150 1410.5650 ;
        RECT 99.3850 1413.8350 99.7150 1414.1650 ;
        RECT 99.3850 1467.8350 99.7150 1468.1650 ;
        RECT 99.3850 1442.6350 99.7150 1442.9650 ;
        RECT 99.3850 1421.0350 99.7150 1421.3650 ;
        RECT 99.3850 1424.6350 99.7150 1424.9650 ;
        RECT 99.3850 1428.2350 99.7150 1428.5650 ;
        RECT 99.3850 1431.8350 99.7150 1432.1650 ;
        RECT 99.3850 1435.4350 99.7150 1435.7650 ;
        RECT 99.3850 1439.0350 99.7150 1439.3650 ;
        RECT 99.3850 1446.2350 99.7150 1446.5650 ;
        RECT 99.3850 1449.8350 99.7150 1450.1650 ;
        RECT 99.3850 1453.4350 99.7150 1453.7650 ;
        RECT 99.3850 1457.0350 99.7150 1457.3650 ;
        RECT 99.3850 1460.6350 99.7150 1460.9650 ;
        RECT 99.3850 1464.2350 99.7150 1464.5650 ;
        RECT 99.3850 1471.4350 99.7150 1471.7650 ;
        RECT 99.3850 1475.0350 99.7150 1475.3650 ;
        RECT 99.3850 1478.6350 99.7150 1478.9650 ;
        RECT 99.3850 1482.2350 99.7150 1482.5650 ;
        RECT 99.3850 1485.8350 99.7150 1486.1650 ;
        RECT 99.3850 1489.4350 99.7150 1489.7650 ;
        RECT 99.3850 1493.0350 99.7150 1493.3650 ;
        RECT 99.3850 1496.6350 99.7150 1496.9650 ;
        RECT 99.3850 1500.2350 99.7150 1500.5650 ;
        RECT 99.3850 1503.8350 99.7150 1504.1650 ;
        RECT 99.3850 1507.4350 99.7150 1507.7650 ;
        RECT 99.3850 1511.0350 99.7150 1511.3650 ;
        RECT 99.3850 1514.6350 99.7150 1514.9650 ;
        RECT 99.3850 1518.2350 99.7150 1518.5650 ;
        RECT 920.1200 816.2350 920.4500 816.5650 ;
        RECT 920.1200 812.6350 920.4500 812.9650 ;
        RECT 920.1200 819.8350 920.4500 820.1650 ;
        RECT 920.1200 823.4350 920.4500 823.7650 ;
        RECT 920.1200 827.0350 920.4500 827.3650 ;
        RECT 920.1200 830.6350 920.4500 830.9650 ;
        RECT 920.1200 834.2350 920.4500 834.5650 ;
        RECT 920.1200 841.4350 920.4500 841.7650 ;
        RECT 920.1200 837.8350 920.4500 838.1650 ;
        RECT 920.1200 845.0350 920.4500 845.3650 ;
        RECT 920.1200 848.6350 920.4500 848.9650 ;
        RECT 920.1200 852.2350 920.4500 852.5650 ;
        RECT 920.1200 855.8350 920.4500 856.1650 ;
        RECT 920.1200 859.4350 920.4500 859.7650 ;
        RECT 920.1200 866.6350 920.4500 866.9650 ;
        RECT 920.1200 863.0350 920.4500 863.3650 ;
        RECT 920.1200 870.2350 920.4500 870.5650 ;
        RECT 920.1200 873.8350 920.4500 874.1650 ;
        RECT 920.1200 877.4350 920.4500 877.7650 ;
        RECT 920.1200 881.0350 920.4500 881.3650 ;
        RECT 920.1200 884.6350 920.4500 884.9650 ;
        RECT 920.1200 888.2350 920.4500 888.5650 ;
        RECT 920.1200 891.8350 920.4500 892.1650 ;
        RECT 920.1200 895.4350 920.4500 895.7650 ;
        RECT 920.1200 899.0350 920.4500 899.3650 ;
        RECT 920.1200 902.6350 920.4500 902.9650 ;
        RECT 920.1200 906.2350 920.4500 906.5650 ;
        RECT 920.1200 909.8350 920.4500 910.1650 ;
        RECT 920.1200 913.4350 920.4500 913.7650 ;
        RECT 920.1200 917.0350 920.4500 917.3650 ;
        RECT 920.1200 920.6350 920.4500 920.9650 ;
        RECT 920.1200 924.2350 920.4500 924.5650 ;
        RECT 920.1200 927.8350 920.4500 928.1650 ;
        RECT 920.1200 931.4350 920.4500 931.7650 ;
        RECT 920.1200 935.0350 920.4500 935.3650 ;
        RECT 920.1200 938.6350 920.4500 938.9650 ;
        RECT 920.1200 942.2350 920.4500 942.5650 ;
        RECT 920.1200 945.8350 920.4500 946.1650 ;
        RECT 920.1200 949.4350 920.4500 949.7650 ;
        RECT 920.1200 953.0350 920.4500 953.3650 ;
        RECT 920.1200 956.6350 920.4500 956.9650 ;
        RECT 920.1200 960.2350 920.4500 960.5650 ;
        RECT 920.1200 963.8350 920.4500 964.1650 ;
        RECT 920.1200 967.4350 920.4500 967.7650 ;
        RECT 920.1200 971.0350 920.4500 971.3650 ;
        RECT 920.1200 974.6350 920.4500 974.9650 ;
        RECT 920.1200 978.2350 920.4500 978.5650 ;
        RECT 920.1200 981.8350 920.4500 982.1650 ;
        RECT 920.1200 985.4350 920.4500 985.7650 ;
        RECT 920.1200 999.8350 920.4500 1000.1650 ;
        RECT 920.1200 989.0350 920.4500 989.3650 ;
        RECT 920.1200 992.6350 920.4500 992.9650 ;
        RECT 920.1200 996.2350 920.4500 996.5650 ;
        RECT 920.1200 1003.4350 920.4500 1003.7650 ;
        RECT 920.1200 1007.0350 920.4500 1007.3650 ;
        RECT 920.1200 1010.6350 920.4500 1010.9650 ;
        RECT 920.1200 1014.2350 920.4500 1014.5650 ;
        RECT 920.1200 1017.8350 920.4500 1018.1650 ;
        RECT 920.1200 1100.6350 920.4500 1100.9650 ;
        RECT 920.1200 1104.2350 920.4500 1104.5650 ;
        RECT 920.1200 1107.8350 920.4500 1108.1650 ;
        RECT 920.1200 1111.4350 920.4500 1111.7650 ;
        RECT 920.1200 1115.0350 920.4500 1115.3650 ;
        RECT 920.1200 1118.6350 920.4500 1118.9650 ;
        RECT 920.1200 1122.2350 920.4500 1122.5650 ;
        RECT 920.1200 1125.8350 920.4500 1126.1650 ;
        RECT 920.1200 1129.4350 920.4500 1129.7650 ;
        RECT 920.1200 1133.0350 920.4500 1133.3650 ;
        RECT 920.1200 1136.6350 920.4500 1136.9650 ;
        RECT 920.1200 1140.2350 920.4500 1140.5650 ;
        RECT 920.1200 1143.8350 920.4500 1144.1650 ;
        RECT 920.1200 1147.4350 920.4500 1147.7650 ;
        RECT 920.1200 1151.0350 920.4500 1151.3650 ;
        RECT 920.1200 1154.6350 920.4500 1154.9650 ;
        RECT 920.1200 1158.2350 920.4500 1158.5650 ;
        RECT 920.1200 1161.8350 920.4500 1162.1650 ;
        RECT 920.1200 1165.4350 920.4500 1165.7650 ;
        RECT 920.1200 1169.0350 920.4500 1169.3650 ;
        RECT 920.1200 1172.6350 920.4500 1172.9650 ;
        RECT 920.1200 1176.2350 920.4500 1176.5650 ;
        RECT 920.1200 1179.8350 920.4500 1180.1650 ;
        RECT 920.1200 1183.4350 920.4500 1183.7650 ;
        RECT 920.1200 1187.0350 920.4500 1187.3650 ;
        RECT 920.1200 1190.6350 920.4500 1190.9650 ;
        RECT 920.1200 1194.2350 920.4500 1194.5650 ;
        RECT 920.1200 1197.8350 920.4500 1198.1650 ;
        RECT 920.1200 1201.4350 920.4500 1201.7650 ;
        RECT 920.1200 1208.6350 920.4500 1208.9650 ;
        RECT 920.1200 1205.0350 920.4500 1205.3650 ;
        RECT 920.1200 1212.2350 920.4500 1212.5650 ;
        RECT 920.1200 1417.4350 920.4500 1417.7650 ;
        RECT 920.1200 1215.8350 920.4500 1216.1650 ;
        RECT 920.1200 1219.4350 920.4500 1219.7650 ;
        RECT 920.1200 1223.0350 920.4500 1223.3650 ;
        RECT 920.1200 1226.6350 920.4500 1226.9650 ;
        RECT 920.1200 1233.8350 920.4500 1234.1650 ;
        RECT 920.1200 1230.2350 920.4500 1230.5650 ;
        RECT 920.1200 1237.4350 920.4500 1237.7650 ;
        RECT 920.1200 1241.0350 920.4500 1241.3650 ;
        RECT 920.1200 1244.6350 920.4500 1244.9650 ;
        RECT 920.1200 1248.2350 920.4500 1248.5650 ;
        RECT 920.1200 1251.8350 920.4500 1252.1650 ;
        RECT 920.1200 1259.0350 920.4500 1259.3650 ;
        RECT 920.1200 1255.4350 920.4500 1255.7650 ;
        RECT 920.1200 1262.6350 920.4500 1262.9650 ;
        RECT 920.1200 1266.2350 920.4500 1266.5650 ;
        RECT 920.1200 1269.8350 920.4500 1270.1650 ;
        RECT 920.1200 1273.4350 920.4500 1273.7650 ;
        RECT 920.1200 1277.0350 920.4500 1277.3650 ;
        RECT 920.1200 1280.6350 920.4500 1280.9650 ;
        RECT 920.1200 1284.2350 920.4500 1284.5650 ;
        RECT 920.1200 1287.8350 920.4500 1288.1650 ;
        RECT 920.1200 1291.4350 920.4500 1291.7650 ;
        RECT 920.1200 1295.0350 920.4500 1295.3650 ;
        RECT 920.1200 1298.6350 920.4500 1298.9650 ;
        RECT 920.1200 1302.2350 920.4500 1302.5650 ;
        RECT 920.1200 1305.8350 920.4500 1306.1650 ;
        RECT 920.1200 1309.4350 920.4500 1309.7650 ;
        RECT 920.1200 1313.0350 920.4500 1313.3650 ;
        RECT 920.1200 1316.6350 920.4500 1316.9650 ;
        RECT 920.1200 1320.2350 920.4500 1320.5650 ;
        RECT 920.1200 1323.8350 920.4500 1324.1650 ;
        RECT 920.1200 1327.4350 920.4500 1327.7650 ;
        RECT 920.1200 1331.0350 920.4500 1331.3650 ;
        RECT 920.1200 1334.6350 920.4500 1334.9650 ;
        RECT 920.1200 1338.2350 920.4500 1338.5650 ;
        RECT 920.1200 1341.8350 920.4500 1342.1650 ;
        RECT 920.1200 1345.4350 920.4500 1345.7650 ;
        RECT 920.1200 1349.0350 920.4500 1349.3650 ;
        RECT 920.1200 1352.6350 920.4500 1352.9650 ;
        RECT 920.1200 1356.2350 920.4500 1356.5650 ;
        RECT 920.1200 1359.8350 920.4500 1360.1650 ;
        RECT 920.1200 1363.4350 920.4500 1363.7650 ;
        RECT 920.1200 1367.0350 920.4500 1367.3650 ;
        RECT 920.1200 1370.6350 920.4500 1370.9650 ;
        RECT 920.1200 1374.2350 920.4500 1374.5650 ;
        RECT 920.1200 1377.8350 920.4500 1378.1650 ;
        RECT 920.1200 1381.4350 920.4500 1381.7650 ;
        RECT 920.1200 1385.0350 920.4500 1385.3650 ;
        RECT 920.1200 1388.6350 920.4500 1388.9650 ;
        RECT 920.1200 1392.2350 920.4500 1392.5650 ;
        RECT 920.1200 1395.8350 920.4500 1396.1650 ;
        RECT 920.1200 1399.4350 920.4500 1399.7650 ;
        RECT 920.1200 1403.0350 920.4500 1403.3650 ;
        RECT 920.1200 1406.6350 920.4500 1406.9650 ;
        RECT 920.1200 1410.2350 920.4500 1410.5650 ;
        RECT 920.1200 1413.8350 920.4500 1414.1650 ;
        RECT 920.1200 1467.8350 920.4500 1468.1650 ;
        RECT 920.1200 1442.6350 920.4500 1442.9650 ;
        RECT 920.1200 1421.0350 920.4500 1421.3650 ;
        RECT 920.1200 1424.6350 920.4500 1424.9650 ;
        RECT 920.1200 1428.2350 920.4500 1428.5650 ;
        RECT 920.1200 1431.8350 920.4500 1432.1650 ;
        RECT 920.1200 1435.4350 920.4500 1435.7650 ;
        RECT 920.1200 1439.0350 920.4500 1439.3650 ;
        RECT 920.1200 1446.2350 920.4500 1446.5650 ;
        RECT 920.1200 1449.8350 920.4500 1450.1650 ;
        RECT 920.1200 1453.4350 920.4500 1453.7650 ;
        RECT 920.1200 1457.0350 920.4500 1457.3650 ;
        RECT 920.1200 1460.6350 920.4500 1460.9650 ;
        RECT 920.1200 1464.2350 920.4500 1464.5650 ;
        RECT 920.1200 1471.4350 920.4500 1471.7650 ;
        RECT 920.1200 1475.0350 920.4500 1475.3650 ;
        RECT 920.1200 1478.6350 920.4500 1478.9650 ;
        RECT 920.1200 1482.2350 920.4500 1482.5650 ;
        RECT 920.1200 1485.8350 920.4500 1486.1650 ;
        RECT 920.1200 1489.4350 920.4500 1489.7650 ;
        RECT 920.1200 1493.0350 920.4500 1493.3650 ;
        RECT 920.1200 1496.6350 920.4500 1496.9650 ;
        RECT 920.1200 1500.2350 920.4500 1500.5650 ;
        RECT 920.1200 1503.8350 920.4500 1504.1650 ;
        RECT 920.1200 1507.4350 920.4500 1507.7650 ;
        RECT 920.1200 1511.0350 920.4500 1511.3650 ;
        RECT 920.1200 1514.6350 920.4500 1514.9650 ;
        RECT 920.1200 1518.2350 920.4500 1518.5650 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 908.9850 609.8350 909.9850 610.1650 ;
        RECT 795.1300 609.8350 796.1300 610.1650 ;
        RECT 681.2750 609.8350 682.2750 610.1650 ;
        RECT 567.4200 609.8350 568.4200 610.1650 ;
        RECT 453.5650 609.8350 454.5650 610.1650 ;
        RECT 339.7100 609.8350 340.7100 610.1650 ;
        RECT 225.8550 609.8350 226.8550 610.1650 ;
        RECT 112.0000 609.8350 113.0000 610.1650 ;
        RECT 112.0000 610.0000 113.0000 1010.0000 ;
        RECT 225.8550 610.0000 226.8550 1010.0000 ;
        RECT 339.7100 610.0000 340.7100 1010.0000 ;
        RECT 453.5650 610.0000 454.5650 1010.0000 ;
        RECT 567.4200 610.0000 568.4200 1010.0000 ;
        RECT 681.2750 610.0000 682.2750 1010.0000 ;
        RECT 795.1300 610.0000 796.1300 1010.0000 ;
        RECT 908.9850 610.0000 909.9850 1010.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 908.9850 1109.8350 909.9850 1110.1650 ;
        RECT 795.1300 1109.8350 796.1300 1110.1650 ;
        RECT 681.2750 1109.8350 682.2750 1110.1650 ;
        RECT 567.4200 1109.8350 568.4200 1110.1650 ;
        RECT 453.5650 1109.8350 454.5650 1110.1650 ;
        RECT 339.7100 1109.8350 340.7100 1110.1650 ;
        RECT 225.8550 1109.8350 226.8550 1110.1650 ;
        RECT 112.0000 1109.8350 113.0000 1110.1650 ;
        RECT 112.0000 1110.0000 113.0000 1510.0000 ;
        RECT 225.8550 1110.0000 226.8550 1510.0000 ;
        RECT 339.7100 1110.0000 340.7100 1510.0000 ;
        RECT 453.5650 1110.0000 454.5650 1510.0000 ;
        RECT 567.4200 1110.0000 568.4200 1510.0000 ;
        RECT 681.2750 1110.0000 682.2750 1510.0000 ;
        RECT 795.1300 1110.0000 796.1300 1510.0000 ;
        RECT 908.9850 1110.0000 909.9850 1510.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'


# P/G pin shape extracted from block 'sram_w16'
    PORT
      LAYER M4 ;
        RECT 908.9850 109.8350 909.9850 110.1650 ;
        RECT 795.1300 109.8350 796.1300 110.1650 ;
        RECT 681.2750 109.8350 682.2750 110.1650 ;
        RECT 567.4200 109.8350 568.4200 110.1650 ;
        RECT 453.5650 109.8350 454.5650 110.1650 ;
        RECT 339.7100 109.8350 340.7100 110.1650 ;
        RECT 225.8550 109.8350 226.8550 110.1650 ;
        RECT 112.0000 109.8350 113.0000 110.1650 ;
        RECT 112.0000 110.0000 113.0000 510.0000 ;
        RECT 225.8550 110.0000 226.8550 510.0000 ;
        RECT 339.7100 110.0000 340.7100 510.0000 ;
        RECT 453.5650 110.0000 454.5650 510.0000 ;
        RECT 567.4200 110.0000 568.4200 510.0000 ;
        RECT 681.2750 110.0000 682.2750 510.0000 ;
        RECT 795.1300 110.0000 796.1300 510.0000 ;
        RECT 908.9850 110.0000 909.9850 510.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16'

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1020.0000 1620.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1020.0000 1620.0000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1020.0000 1620.0000 ;
    LAYER M4 ;
      RECT 0.0000 1610.5000 1020.0000 1620.0000 ;
      RECT 900.5000 1520.4850 999.5000 1610.5000 ;
      RECT 20.5000 1520.4850 119.5000 1610.5000 ;
      RECT 920.5450 1519.9150 999.5000 1520.4850 ;
      RECT 900.5000 1519.9150 919.9750 1520.4850 ;
      RECT 99.8600 1519.9150 119.5000 1520.4850 ;
      RECT 20.5000 1519.9150 99.2900 1520.4850 ;
      RECT 900.5000 1518.6850 999.5000 1519.9150 ;
      RECT 20.5000 1518.6850 119.5000 1519.9150 ;
      RECT 920.5700 1518.1150 999.5000 1518.6850 ;
      RECT 900.5000 1518.1150 920.0000 1518.6850 ;
      RECT 99.8350 1518.1150 119.5000 1518.6850 ;
      RECT 20.5000 1518.1150 99.2650 1518.6850 ;
      RECT 900.5000 1516.8850 999.5000 1518.1150 ;
      RECT 20.5000 1516.8850 119.5000 1518.1150 ;
      RECT 920.5700 1516.3150 999.5000 1516.8850 ;
      RECT 900.5000 1516.3150 920.0000 1516.8850 ;
      RECT 99.8350 1516.3150 119.5000 1516.8850 ;
      RECT 20.5000 1516.3150 99.2650 1516.8850 ;
      RECT 900.5000 1515.0850 999.5000 1516.3150 ;
      RECT 20.5000 1515.0850 119.5000 1516.3150 ;
      RECT 920.5700 1514.5150 999.5000 1515.0850 ;
      RECT 900.5000 1514.5150 920.0000 1515.0850 ;
      RECT 99.8350 1514.5150 119.5000 1515.0850 ;
      RECT 20.5000 1514.5150 99.2650 1515.0850 ;
      RECT 900.5000 1513.2850 999.5000 1514.5150 ;
      RECT 20.5000 1513.2850 119.5000 1514.5150 ;
      RECT 920.5700 1512.7150 999.5000 1513.2850 ;
      RECT 900.5000 1512.7150 920.0000 1513.2850 ;
      RECT 99.8350 1512.7150 119.5000 1513.2850 ;
      RECT 20.5000 1512.7150 99.2650 1513.2850 ;
      RECT 900.5000 1511.4850 999.5000 1512.7150 ;
      RECT 20.5000 1511.4850 119.5000 1512.7150 ;
      RECT 920.5700 1510.9150 999.5000 1511.4850 ;
      RECT 900.5000 1510.9150 920.0000 1511.4850 ;
      RECT 99.8350 1510.9150 119.5000 1511.4850 ;
      RECT 20.5000 1510.9150 99.2650 1511.4850 ;
      RECT 900.5000 1509.6850 999.5000 1510.9150 ;
      RECT 20.5000 1509.6850 119.5000 1510.9150 ;
      RECT 920.5700 1509.1150 999.5000 1509.6850 ;
      RECT 900.5000 1509.1150 920.0000 1509.6850 ;
      RECT 99.8350 1509.1150 119.5000 1509.6850 ;
      RECT 20.5000 1509.1150 99.2650 1509.6850 ;
      RECT 900.5000 1507.8850 999.5000 1509.1150 ;
      RECT 20.5000 1507.8850 119.5000 1509.1150 ;
      RECT 920.5700 1507.3150 999.5000 1507.8850 ;
      RECT 900.5000 1507.3150 920.0000 1507.8850 ;
      RECT 99.8350 1507.3150 119.5000 1507.8850 ;
      RECT 20.5000 1507.3150 99.2650 1507.8850 ;
      RECT 900.5000 1506.0850 999.5000 1507.3150 ;
      RECT 20.5000 1506.0850 119.5000 1507.3150 ;
      RECT 920.5700 1505.5150 999.5000 1506.0850 ;
      RECT 900.5000 1505.5150 920.0000 1506.0850 ;
      RECT 99.8350 1505.5150 119.5000 1506.0850 ;
      RECT 20.5000 1505.5150 99.2650 1506.0850 ;
      RECT 900.5000 1504.2850 999.5000 1505.5150 ;
      RECT 20.5000 1504.2850 119.5000 1505.5150 ;
      RECT 920.5700 1503.7150 999.5000 1504.2850 ;
      RECT 900.5000 1503.7150 920.0000 1504.2850 ;
      RECT 99.8350 1503.7150 119.5000 1504.2850 ;
      RECT 20.5000 1503.7150 99.2650 1504.2850 ;
      RECT 900.5000 1502.4850 999.5000 1503.7150 ;
      RECT 20.5000 1502.4850 119.5000 1503.7150 ;
      RECT 920.5700 1501.9150 999.5000 1502.4850 ;
      RECT 900.5000 1501.9150 920.0000 1502.4850 ;
      RECT 99.8350 1501.9150 119.5000 1502.4850 ;
      RECT 20.5000 1501.9150 99.2650 1502.4850 ;
      RECT 900.5000 1500.6850 999.5000 1501.9150 ;
      RECT 20.5000 1500.6850 119.5000 1501.9150 ;
      RECT 920.5700 1500.1150 999.5000 1500.6850 ;
      RECT 900.5000 1500.1150 920.0000 1500.6850 ;
      RECT 99.8350 1500.1150 119.5000 1500.6850 ;
      RECT 20.5000 1500.1150 99.2650 1500.6850 ;
      RECT 900.5000 1498.8850 999.5000 1500.1150 ;
      RECT 20.5000 1498.8850 119.5000 1500.1150 ;
      RECT 920.5700 1498.3150 999.5000 1498.8850 ;
      RECT 900.5000 1498.3150 920.0000 1498.8850 ;
      RECT 99.8350 1498.3150 119.5000 1498.8850 ;
      RECT 20.5000 1498.3150 99.2650 1498.8850 ;
      RECT 900.5000 1497.0850 999.5000 1498.3150 ;
      RECT 20.5000 1497.0850 119.5000 1498.3150 ;
      RECT 920.5700 1496.5150 999.5000 1497.0850 ;
      RECT 900.5000 1496.5150 920.0000 1497.0850 ;
      RECT 99.8350 1496.5150 119.5000 1497.0850 ;
      RECT 20.5000 1496.5150 99.2650 1497.0850 ;
      RECT 900.5000 1495.2850 999.5000 1496.5150 ;
      RECT 20.5000 1495.2850 119.5000 1496.5150 ;
      RECT 920.5700 1494.7150 999.5000 1495.2850 ;
      RECT 900.5000 1494.7150 920.0000 1495.2850 ;
      RECT 99.8350 1494.7150 119.5000 1495.2850 ;
      RECT 20.5000 1494.7150 99.2650 1495.2850 ;
      RECT 900.5000 1493.4850 999.5000 1494.7150 ;
      RECT 20.5000 1493.4850 119.5000 1494.7150 ;
      RECT 920.5700 1492.9150 999.5000 1493.4850 ;
      RECT 900.5000 1492.9150 920.0000 1493.4850 ;
      RECT 99.8350 1492.9150 119.5000 1493.4850 ;
      RECT 20.5000 1492.9150 99.2650 1493.4850 ;
      RECT 900.5000 1491.6850 999.5000 1492.9150 ;
      RECT 20.5000 1491.6850 119.5000 1492.9150 ;
      RECT 920.5700 1491.1150 999.5000 1491.6850 ;
      RECT 900.5000 1491.1150 920.0000 1491.6850 ;
      RECT 99.8350 1491.1150 119.5000 1491.6850 ;
      RECT 20.5000 1491.1150 99.2650 1491.6850 ;
      RECT 900.5000 1489.8850 999.5000 1491.1150 ;
      RECT 20.5000 1489.8850 119.5000 1491.1150 ;
      RECT 920.5700 1489.3150 999.5000 1489.8850 ;
      RECT 900.5000 1489.3150 920.0000 1489.8850 ;
      RECT 99.8350 1489.3150 119.5000 1489.8850 ;
      RECT 20.5000 1489.3150 99.2650 1489.8850 ;
      RECT 900.5000 1488.0850 999.5000 1489.3150 ;
      RECT 20.5000 1488.0850 119.5000 1489.3150 ;
      RECT 920.5700 1487.5150 999.5000 1488.0850 ;
      RECT 900.5000 1487.5150 920.0000 1488.0850 ;
      RECT 99.8350 1487.5150 119.5000 1488.0850 ;
      RECT 20.5000 1487.5150 99.2650 1488.0850 ;
      RECT 900.5000 1486.2850 999.5000 1487.5150 ;
      RECT 20.5000 1486.2850 119.5000 1487.5150 ;
      RECT 920.5700 1485.7150 999.5000 1486.2850 ;
      RECT 900.5000 1485.7150 920.0000 1486.2850 ;
      RECT 99.8350 1485.7150 119.5000 1486.2850 ;
      RECT 20.5000 1485.7150 99.2650 1486.2850 ;
      RECT 900.5000 1484.4850 999.5000 1485.7150 ;
      RECT 20.5000 1484.4850 119.5000 1485.7150 ;
      RECT 920.5700 1483.9150 999.5000 1484.4850 ;
      RECT 900.5000 1483.9150 920.0000 1484.4850 ;
      RECT 99.8350 1483.9150 119.5000 1484.4850 ;
      RECT 20.5000 1483.9150 99.2650 1484.4850 ;
      RECT 900.5000 1482.6850 999.5000 1483.9150 ;
      RECT 20.5000 1482.6850 119.5000 1483.9150 ;
      RECT 920.5700 1482.1150 999.5000 1482.6850 ;
      RECT 900.5000 1482.1150 920.0000 1482.6850 ;
      RECT 99.8350 1482.1150 119.5000 1482.6850 ;
      RECT 20.5000 1482.1150 99.2650 1482.6850 ;
      RECT 900.5000 1480.8850 999.5000 1482.1150 ;
      RECT 20.5000 1480.8850 119.5000 1482.1150 ;
      RECT 920.5700 1480.3150 999.5000 1480.8850 ;
      RECT 900.5000 1480.3150 920.0000 1480.8850 ;
      RECT 99.8350 1480.3150 119.5000 1480.8850 ;
      RECT 20.5000 1480.3150 99.2650 1480.8850 ;
      RECT 900.5000 1479.0850 999.5000 1480.3150 ;
      RECT 20.5000 1479.0850 119.5000 1480.3150 ;
      RECT 920.5700 1478.5150 999.5000 1479.0850 ;
      RECT 900.5000 1478.5150 920.0000 1479.0850 ;
      RECT 99.8350 1478.5150 119.5000 1479.0850 ;
      RECT 20.5000 1478.5150 99.2650 1479.0850 ;
      RECT 900.5000 1477.2850 999.5000 1478.5150 ;
      RECT 20.5000 1477.2850 119.5000 1478.5150 ;
      RECT 920.5700 1476.7150 999.5000 1477.2850 ;
      RECT 900.5000 1476.7150 920.0000 1477.2850 ;
      RECT 99.8350 1476.7150 119.5000 1477.2850 ;
      RECT 20.5000 1476.7150 99.2650 1477.2850 ;
      RECT 900.5000 1475.4850 999.5000 1476.7150 ;
      RECT 20.5000 1475.4850 119.5000 1476.7150 ;
      RECT 920.5700 1474.9150 999.5000 1475.4850 ;
      RECT 900.5000 1474.9150 920.0000 1475.4850 ;
      RECT 99.8350 1474.9150 119.5000 1475.4850 ;
      RECT 20.5000 1474.9150 99.2650 1475.4850 ;
      RECT 900.5000 1473.6850 999.5000 1474.9150 ;
      RECT 20.5000 1473.6850 119.5000 1474.9150 ;
      RECT 920.5700 1473.1150 999.5000 1473.6850 ;
      RECT 900.5000 1473.1150 920.0000 1473.6850 ;
      RECT 99.8350 1473.1150 119.5000 1473.6850 ;
      RECT 20.5000 1473.1150 99.2650 1473.6850 ;
      RECT 900.5000 1471.8850 999.5000 1473.1150 ;
      RECT 20.5000 1471.8850 119.5000 1473.1150 ;
      RECT 920.5700 1471.3150 999.5000 1471.8850 ;
      RECT 900.5000 1471.3150 920.0000 1471.8850 ;
      RECT 99.8350 1471.3150 119.5000 1471.8850 ;
      RECT 20.5000 1471.3150 99.2650 1471.8850 ;
      RECT 900.5000 1470.0850 999.5000 1471.3150 ;
      RECT 20.5000 1470.0850 119.5000 1471.3150 ;
      RECT 920.5700 1469.5150 999.5000 1470.0850 ;
      RECT 900.5000 1469.5150 920.0000 1470.0850 ;
      RECT 99.8350 1469.5150 119.5000 1470.0850 ;
      RECT 20.5000 1469.5150 99.2650 1470.0850 ;
      RECT 900.5000 1468.2850 999.5000 1469.5150 ;
      RECT 20.5000 1468.2850 119.5000 1469.5150 ;
      RECT 920.5700 1467.7150 999.5000 1468.2850 ;
      RECT 900.5000 1467.7150 920.0000 1468.2850 ;
      RECT 99.8350 1467.7150 119.5000 1468.2850 ;
      RECT 20.5000 1467.7150 99.2650 1468.2850 ;
      RECT 900.5000 1466.4850 999.5000 1467.7150 ;
      RECT 20.5000 1466.4850 119.5000 1467.7150 ;
      RECT 920.5700 1465.9150 999.5000 1466.4850 ;
      RECT 900.5000 1465.9150 920.0000 1466.4850 ;
      RECT 99.8350 1465.9150 119.5000 1466.4850 ;
      RECT 20.5000 1465.9150 99.2650 1466.4850 ;
      RECT 900.5000 1464.6850 999.5000 1465.9150 ;
      RECT 20.5000 1464.6850 119.5000 1465.9150 ;
      RECT 920.5700 1464.1150 999.5000 1464.6850 ;
      RECT 900.5000 1464.1150 920.0000 1464.6850 ;
      RECT 99.8350 1464.1150 119.5000 1464.6850 ;
      RECT 20.5000 1464.1150 99.2650 1464.6850 ;
      RECT 900.5000 1462.8850 999.5000 1464.1150 ;
      RECT 20.5000 1462.8850 119.5000 1464.1150 ;
      RECT 920.5700 1462.3150 999.5000 1462.8850 ;
      RECT 900.5000 1462.3150 920.0000 1462.8850 ;
      RECT 99.8350 1462.3150 119.5000 1462.8850 ;
      RECT 20.5000 1462.3150 99.2650 1462.8850 ;
      RECT 900.5000 1461.0850 999.5000 1462.3150 ;
      RECT 20.5000 1461.0850 119.5000 1462.3150 ;
      RECT 920.5700 1460.5150 999.5000 1461.0850 ;
      RECT 900.5000 1460.5150 920.0000 1461.0850 ;
      RECT 99.8350 1460.5150 119.5000 1461.0850 ;
      RECT 20.5000 1460.5150 99.2650 1461.0850 ;
      RECT 900.5000 1459.2850 999.5000 1460.5150 ;
      RECT 20.5000 1459.2850 119.5000 1460.5150 ;
      RECT 920.5700 1458.7150 999.5000 1459.2850 ;
      RECT 900.5000 1458.7150 920.0000 1459.2850 ;
      RECT 99.8350 1458.7150 119.5000 1459.2850 ;
      RECT 20.5000 1458.7150 99.2650 1459.2850 ;
      RECT 900.5000 1457.4850 999.5000 1458.7150 ;
      RECT 20.5000 1457.4850 119.5000 1458.7150 ;
      RECT 920.5700 1456.9150 999.5000 1457.4850 ;
      RECT 900.5000 1456.9150 920.0000 1457.4850 ;
      RECT 99.8350 1456.9150 119.5000 1457.4850 ;
      RECT 20.5000 1456.9150 99.2650 1457.4850 ;
      RECT 900.5000 1455.6850 999.5000 1456.9150 ;
      RECT 20.5000 1455.6850 119.5000 1456.9150 ;
      RECT 920.5700 1455.1150 999.5000 1455.6850 ;
      RECT 900.5000 1455.1150 920.0000 1455.6850 ;
      RECT 99.8350 1455.1150 119.5000 1455.6850 ;
      RECT 20.5000 1455.1150 99.2650 1455.6850 ;
      RECT 900.5000 1453.8850 999.5000 1455.1150 ;
      RECT 20.5000 1453.8850 119.5000 1455.1150 ;
      RECT 920.5700 1453.3150 999.5000 1453.8850 ;
      RECT 900.5000 1453.3150 920.0000 1453.8850 ;
      RECT 99.8350 1453.3150 119.5000 1453.8850 ;
      RECT 20.5000 1453.3150 99.2650 1453.8850 ;
      RECT 900.5000 1452.0850 999.5000 1453.3150 ;
      RECT 20.5000 1452.0850 119.5000 1453.3150 ;
      RECT 920.5700 1451.5150 999.5000 1452.0850 ;
      RECT 900.5000 1451.5150 920.0000 1452.0850 ;
      RECT 99.8350 1451.5150 119.5000 1452.0850 ;
      RECT 20.5000 1451.5150 99.2650 1452.0850 ;
      RECT 900.5000 1450.2850 999.5000 1451.5150 ;
      RECT 20.5000 1450.2850 119.5000 1451.5150 ;
      RECT 920.5700 1449.7150 999.5000 1450.2850 ;
      RECT 900.5000 1449.7150 920.0000 1450.2850 ;
      RECT 99.8350 1449.7150 119.5000 1450.2850 ;
      RECT 20.5000 1449.7150 99.2650 1450.2850 ;
      RECT 900.5000 1448.4850 999.5000 1449.7150 ;
      RECT 20.5000 1448.4850 119.5000 1449.7150 ;
      RECT 920.5700 1447.9150 999.5000 1448.4850 ;
      RECT 900.5000 1447.9150 920.0000 1448.4850 ;
      RECT 99.8350 1447.9150 119.5000 1448.4850 ;
      RECT 20.5000 1447.9150 99.2650 1448.4850 ;
      RECT 900.5000 1446.6850 999.5000 1447.9150 ;
      RECT 20.5000 1446.6850 119.5000 1447.9150 ;
      RECT 920.5700 1446.1150 999.5000 1446.6850 ;
      RECT 900.5000 1446.1150 920.0000 1446.6850 ;
      RECT 99.8350 1446.1150 119.5000 1446.6850 ;
      RECT 20.5000 1446.1150 99.2650 1446.6850 ;
      RECT 900.5000 1444.8850 999.5000 1446.1150 ;
      RECT 20.5000 1444.8850 119.5000 1446.1150 ;
      RECT 920.5700 1444.3150 999.5000 1444.8850 ;
      RECT 900.5000 1444.3150 920.0000 1444.8850 ;
      RECT 99.8350 1444.3150 119.5000 1444.8850 ;
      RECT 20.5000 1444.3150 99.2650 1444.8850 ;
      RECT 900.5000 1443.0850 999.5000 1444.3150 ;
      RECT 20.5000 1443.0850 119.5000 1444.3150 ;
      RECT 920.5700 1442.5150 999.5000 1443.0850 ;
      RECT 900.5000 1442.5150 920.0000 1443.0850 ;
      RECT 99.8350 1442.5150 119.5000 1443.0850 ;
      RECT 20.5000 1442.5150 99.2650 1443.0850 ;
      RECT 900.5000 1441.2850 999.5000 1442.5150 ;
      RECT 20.5000 1441.2850 119.5000 1442.5150 ;
      RECT 920.5700 1440.7150 999.5000 1441.2850 ;
      RECT 900.5000 1440.7150 920.0000 1441.2850 ;
      RECT 99.8350 1440.7150 119.5000 1441.2850 ;
      RECT 20.5000 1440.7150 99.2650 1441.2850 ;
      RECT 900.5000 1439.4850 999.5000 1440.7150 ;
      RECT 20.5000 1439.4850 119.5000 1440.7150 ;
      RECT 920.5700 1438.9150 999.5000 1439.4850 ;
      RECT 900.5000 1438.9150 920.0000 1439.4850 ;
      RECT 99.8350 1438.9150 119.5000 1439.4850 ;
      RECT 20.5000 1438.9150 99.2650 1439.4850 ;
      RECT 900.5000 1437.6850 999.5000 1438.9150 ;
      RECT 20.5000 1437.6850 119.5000 1438.9150 ;
      RECT 920.5700 1437.1150 999.5000 1437.6850 ;
      RECT 900.5000 1437.1150 920.0000 1437.6850 ;
      RECT 99.8350 1437.1150 119.5000 1437.6850 ;
      RECT 20.5000 1437.1150 99.2650 1437.6850 ;
      RECT 900.5000 1435.8850 999.5000 1437.1150 ;
      RECT 20.5000 1435.8850 119.5000 1437.1150 ;
      RECT 920.5700 1435.3150 999.5000 1435.8850 ;
      RECT 900.5000 1435.3150 920.0000 1435.8850 ;
      RECT 99.8350 1435.3150 119.5000 1435.8850 ;
      RECT 20.5000 1435.3150 99.2650 1435.8850 ;
      RECT 900.5000 1434.0850 999.5000 1435.3150 ;
      RECT 20.5000 1434.0850 119.5000 1435.3150 ;
      RECT 920.5700 1433.5150 999.5000 1434.0850 ;
      RECT 900.5000 1433.5150 920.0000 1434.0850 ;
      RECT 99.8350 1433.5150 119.5000 1434.0850 ;
      RECT 20.5000 1433.5150 99.2650 1434.0850 ;
      RECT 900.5000 1432.2850 999.5000 1433.5150 ;
      RECT 20.5000 1432.2850 119.5000 1433.5150 ;
      RECT 920.5700 1431.7150 999.5000 1432.2850 ;
      RECT 900.5000 1431.7150 920.0000 1432.2850 ;
      RECT 99.8350 1431.7150 119.5000 1432.2850 ;
      RECT 20.5000 1431.7150 99.2650 1432.2850 ;
      RECT 900.5000 1430.4850 999.5000 1431.7150 ;
      RECT 20.5000 1430.4850 119.5000 1431.7150 ;
      RECT 920.5700 1429.9150 999.5000 1430.4850 ;
      RECT 900.5000 1429.9150 920.0000 1430.4850 ;
      RECT 99.8350 1429.9150 119.5000 1430.4850 ;
      RECT 20.5000 1429.9150 99.2650 1430.4850 ;
      RECT 900.5000 1428.6850 999.5000 1429.9150 ;
      RECT 20.5000 1428.6850 119.5000 1429.9150 ;
      RECT 920.5700 1428.1150 999.5000 1428.6850 ;
      RECT 900.5000 1428.1150 920.0000 1428.6850 ;
      RECT 99.8350 1428.1150 119.5000 1428.6850 ;
      RECT 20.5000 1428.1150 99.2650 1428.6850 ;
      RECT 900.5000 1426.8850 999.5000 1428.1150 ;
      RECT 20.5000 1426.8850 119.5000 1428.1150 ;
      RECT 920.5700 1426.3150 999.5000 1426.8850 ;
      RECT 900.5000 1426.3150 920.0000 1426.8850 ;
      RECT 99.8350 1426.3150 119.5000 1426.8850 ;
      RECT 20.5000 1426.3150 99.2650 1426.8850 ;
      RECT 900.5000 1425.0850 999.5000 1426.3150 ;
      RECT 20.5000 1425.0850 119.5000 1426.3150 ;
      RECT 920.5700 1424.5150 999.5000 1425.0850 ;
      RECT 900.5000 1424.5150 920.0000 1425.0850 ;
      RECT 99.8350 1424.5150 119.5000 1425.0850 ;
      RECT 20.5000 1424.5150 99.2650 1425.0850 ;
      RECT 900.5000 1423.2850 999.5000 1424.5150 ;
      RECT 20.5000 1423.2850 119.5000 1424.5150 ;
      RECT 920.5700 1422.7150 999.5000 1423.2850 ;
      RECT 900.5000 1422.7150 920.0000 1423.2850 ;
      RECT 99.8350 1422.7150 119.5000 1423.2850 ;
      RECT 20.5000 1422.7150 99.2650 1423.2850 ;
      RECT 900.5000 1421.4850 999.5000 1422.7150 ;
      RECT 20.5000 1421.4850 119.5000 1422.7150 ;
      RECT 920.5700 1420.9150 999.5000 1421.4850 ;
      RECT 900.5000 1420.9150 920.0000 1421.4850 ;
      RECT 99.8350 1420.9150 119.5000 1421.4850 ;
      RECT 20.5000 1420.9150 99.2650 1421.4850 ;
      RECT 900.5000 1419.6850 999.5000 1420.9150 ;
      RECT 20.5000 1419.6850 119.5000 1420.9150 ;
      RECT 920.5700 1419.1150 999.5000 1419.6850 ;
      RECT 900.5000 1419.1150 920.0000 1419.6850 ;
      RECT 99.8350 1419.1150 119.5000 1419.6850 ;
      RECT 20.5000 1419.1150 99.2650 1419.6850 ;
      RECT 900.5000 1417.8850 999.5000 1419.1150 ;
      RECT 20.5000 1417.8850 119.5000 1419.1150 ;
      RECT 920.5700 1417.3150 999.5000 1417.8850 ;
      RECT 900.5000 1417.3150 920.0000 1417.8850 ;
      RECT 99.8350 1417.3150 119.5000 1417.8850 ;
      RECT 20.5000 1417.3150 99.2650 1417.8850 ;
      RECT 900.5000 1416.0850 999.5000 1417.3150 ;
      RECT 20.5000 1416.0850 119.5000 1417.3150 ;
      RECT 920.5700 1415.5150 999.5000 1416.0850 ;
      RECT 900.5000 1415.5150 920.0000 1416.0850 ;
      RECT 99.8350 1415.5150 119.5000 1416.0850 ;
      RECT 20.5000 1415.5150 99.2650 1416.0850 ;
      RECT 900.5000 1414.2850 999.5000 1415.5150 ;
      RECT 20.5000 1414.2850 119.5000 1415.5150 ;
      RECT 920.5700 1413.7150 999.5000 1414.2850 ;
      RECT 900.5000 1413.7150 920.0000 1414.2850 ;
      RECT 99.8350 1413.7150 119.5000 1414.2850 ;
      RECT 20.5000 1413.7150 99.2650 1414.2850 ;
      RECT 900.5000 1412.4850 999.5000 1413.7150 ;
      RECT 20.5000 1412.4850 119.5000 1413.7150 ;
      RECT 920.5700 1411.9150 999.5000 1412.4850 ;
      RECT 900.5000 1411.9150 920.0000 1412.4850 ;
      RECT 99.8350 1411.9150 119.5000 1412.4850 ;
      RECT 20.5000 1411.9150 99.2650 1412.4850 ;
      RECT 900.5000 1410.6850 999.5000 1411.9150 ;
      RECT 20.5000 1410.6850 119.5000 1411.9150 ;
      RECT 920.5700 1410.1150 999.5000 1410.6850 ;
      RECT 900.5000 1410.1150 920.0000 1410.6850 ;
      RECT 99.8350 1410.1150 119.5000 1410.6850 ;
      RECT 20.5000 1410.1150 99.2650 1410.6850 ;
      RECT 900.5000 1408.8850 999.5000 1410.1150 ;
      RECT 20.5000 1408.8850 119.5000 1410.1150 ;
      RECT 920.5700 1408.3150 999.5000 1408.8850 ;
      RECT 900.5000 1408.3150 920.0000 1408.8850 ;
      RECT 99.8350 1408.3150 119.5000 1408.8850 ;
      RECT 20.5000 1408.3150 99.2650 1408.8850 ;
      RECT 900.5000 1407.0850 999.5000 1408.3150 ;
      RECT 20.5000 1407.0850 119.5000 1408.3150 ;
      RECT 920.5700 1406.5150 999.5000 1407.0850 ;
      RECT 900.5000 1406.5150 920.0000 1407.0850 ;
      RECT 99.8350 1406.5150 119.5000 1407.0850 ;
      RECT 20.5000 1406.5150 99.2650 1407.0850 ;
      RECT 900.5000 1405.2850 999.5000 1406.5150 ;
      RECT 20.5000 1405.2850 119.5000 1406.5150 ;
      RECT 920.5700 1404.7150 999.5000 1405.2850 ;
      RECT 900.5000 1404.7150 920.0000 1405.2850 ;
      RECT 99.8350 1404.7150 119.5000 1405.2850 ;
      RECT 20.5000 1404.7150 99.2650 1405.2850 ;
      RECT 900.5000 1403.4850 999.5000 1404.7150 ;
      RECT 20.5000 1403.4850 119.5000 1404.7150 ;
      RECT 920.5700 1402.9150 999.5000 1403.4850 ;
      RECT 900.5000 1402.9150 920.0000 1403.4850 ;
      RECT 99.8350 1402.9150 119.5000 1403.4850 ;
      RECT 20.5000 1402.9150 99.2650 1403.4850 ;
      RECT 900.5000 1401.6850 999.5000 1402.9150 ;
      RECT 20.5000 1401.6850 119.5000 1402.9150 ;
      RECT 920.5700 1401.1150 999.5000 1401.6850 ;
      RECT 900.5000 1401.1150 920.0000 1401.6850 ;
      RECT 99.8350 1401.1150 119.5000 1401.6850 ;
      RECT 20.5000 1401.1150 99.2650 1401.6850 ;
      RECT 900.5000 1399.8850 999.5000 1401.1150 ;
      RECT 20.5000 1399.8850 119.5000 1401.1150 ;
      RECT 920.5700 1399.3150 999.5000 1399.8850 ;
      RECT 900.5000 1399.3150 920.0000 1399.8850 ;
      RECT 99.8350 1399.3150 119.5000 1399.8850 ;
      RECT 20.5000 1399.3150 99.2650 1399.8850 ;
      RECT 900.5000 1398.0850 999.5000 1399.3150 ;
      RECT 20.5000 1398.0850 119.5000 1399.3150 ;
      RECT 920.5700 1397.5150 999.5000 1398.0850 ;
      RECT 900.5000 1397.5150 920.0000 1398.0850 ;
      RECT 99.8350 1397.5150 119.5000 1398.0850 ;
      RECT 20.5000 1397.5150 99.2650 1398.0850 ;
      RECT 900.5000 1396.2850 999.5000 1397.5150 ;
      RECT 20.5000 1396.2850 119.5000 1397.5150 ;
      RECT 920.5700 1395.7150 999.5000 1396.2850 ;
      RECT 900.5000 1395.7150 920.0000 1396.2850 ;
      RECT 99.8350 1395.7150 119.5000 1396.2850 ;
      RECT 20.5000 1395.7150 99.2650 1396.2850 ;
      RECT 900.5000 1394.4850 999.5000 1395.7150 ;
      RECT 20.5000 1394.4850 119.5000 1395.7150 ;
      RECT 920.5700 1393.9150 999.5000 1394.4850 ;
      RECT 900.5000 1393.9150 920.0000 1394.4850 ;
      RECT 99.8350 1393.9150 119.5000 1394.4850 ;
      RECT 20.5000 1393.9150 99.2650 1394.4850 ;
      RECT 900.5000 1392.6850 999.5000 1393.9150 ;
      RECT 20.5000 1392.6850 119.5000 1393.9150 ;
      RECT 920.5700 1392.1150 999.5000 1392.6850 ;
      RECT 900.5000 1392.1150 920.0000 1392.6850 ;
      RECT 99.8350 1392.1150 119.5000 1392.6850 ;
      RECT 20.5000 1392.1150 99.2650 1392.6850 ;
      RECT 900.5000 1390.8850 999.5000 1392.1150 ;
      RECT 20.5000 1390.8850 119.5000 1392.1150 ;
      RECT 920.5700 1390.3150 999.5000 1390.8850 ;
      RECT 900.5000 1390.3150 920.0000 1390.8850 ;
      RECT 99.8350 1390.3150 119.5000 1390.8850 ;
      RECT 20.5000 1390.3150 99.2650 1390.8850 ;
      RECT 900.5000 1389.0850 999.5000 1390.3150 ;
      RECT 20.5000 1389.0850 119.5000 1390.3150 ;
      RECT 920.5700 1388.5150 999.5000 1389.0850 ;
      RECT 900.5000 1388.5150 920.0000 1389.0850 ;
      RECT 99.8350 1388.5150 119.5000 1389.0850 ;
      RECT 20.5000 1388.5150 99.2650 1389.0850 ;
      RECT 900.5000 1387.2850 999.5000 1388.5150 ;
      RECT 20.5000 1387.2850 119.5000 1388.5150 ;
      RECT 920.5700 1386.7150 999.5000 1387.2850 ;
      RECT 900.5000 1386.7150 920.0000 1387.2850 ;
      RECT 99.8350 1386.7150 119.5000 1387.2850 ;
      RECT 20.5000 1386.7150 99.2650 1387.2850 ;
      RECT 900.5000 1385.4850 999.5000 1386.7150 ;
      RECT 20.5000 1385.4850 119.5000 1386.7150 ;
      RECT 920.5700 1384.9150 999.5000 1385.4850 ;
      RECT 900.5000 1384.9150 920.0000 1385.4850 ;
      RECT 99.8350 1384.9150 119.5000 1385.4850 ;
      RECT 20.5000 1384.9150 99.2650 1385.4850 ;
      RECT 900.5000 1383.6850 999.5000 1384.9150 ;
      RECT 20.5000 1383.6850 119.5000 1384.9150 ;
      RECT 920.5700 1383.1150 999.5000 1383.6850 ;
      RECT 900.5000 1383.1150 920.0000 1383.6850 ;
      RECT 99.8350 1383.1150 119.5000 1383.6850 ;
      RECT 20.5000 1383.1150 99.2650 1383.6850 ;
      RECT 900.5000 1381.8850 999.5000 1383.1150 ;
      RECT 20.5000 1381.8850 119.5000 1383.1150 ;
      RECT 920.5700 1381.3150 999.5000 1381.8850 ;
      RECT 900.5000 1381.3150 920.0000 1381.8850 ;
      RECT 99.8350 1381.3150 119.5000 1381.8850 ;
      RECT 20.5000 1381.3150 99.2650 1381.8850 ;
      RECT 900.5000 1380.0850 999.5000 1381.3150 ;
      RECT 20.5000 1380.0850 119.5000 1381.3150 ;
      RECT 920.5700 1379.5150 999.5000 1380.0850 ;
      RECT 900.5000 1379.5150 920.0000 1380.0850 ;
      RECT 99.8350 1379.5150 119.5000 1380.0850 ;
      RECT 20.5000 1379.5150 99.2650 1380.0850 ;
      RECT 900.5000 1378.2850 999.5000 1379.5150 ;
      RECT 20.5000 1378.2850 119.5000 1379.5150 ;
      RECT 920.5700 1377.7150 999.5000 1378.2850 ;
      RECT 900.5000 1377.7150 920.0000 1378.2850 ;
      RECT 99.8350 1377.7150 119.5000 1378.2850 ;
      RECT 20.5000 1377.7150 99.2650 1378.2850 ;
      RECT 900.5000 1376.4850 999.5000 1377.7150 ;
      RECT 20.5000 1376.4850 119.5000 1377.7150 ;
      RECT 920.5700 1375.9150 999.5000 1376.4850 ;
      RECT 900.5000 1375.9150 920.0000 1376.4850 ;
      RECT 99.8350 1375.9150 119.5000 1376.4850 ;
      RECT 20.5000 1375.9150 99.2650 1376.4850 ;
      RECT 900.5000 1374.6850 999.5000 1375.9150 ;
      RECT 20.5000 1374.6850 119.5000 1375.9150 ;
      RECT 920.5700 1374.1150 999.5000 1374.6850 ;
      RECT 900.5000 1374.1150 920.0000 1374.6850 ;
      RECT 99.8350 1374.1150 119.5000 1374.6850 ;
      RECT 20.5000 1374.1150 99.2650 1374.6850 ;
      RECT 900.5000 1372.8850 999.5000 1374.1150 ;
      RECT 20.5000 1372.8850 119.5000 1374.1150 ;
      RECT 920.5700 1372.3150 999.5000 1372.8850 ;
      RECT 900.5000 1372.3150 920.0000 1372.8850 ;
      RECT 99.8350 1372.3150 119.5000 1372.8850 ;
      RECT 20.5000 1372.3150 99.2650 1372.8850 ;
      RECT 900.5000 1371.0850 999.5000 1372.3150 ;
      RECT 20.5000 1371.0850 119.5000 1372.3150 ;
      RECT 920.5700 1370.5150 999.5000 1371.0850 ;
      RECT 900.5000 1370.5150 920.0000 1371.0850 ;
      RECT 99.8350 1370.5150 119.5000 1371.0850 ;
      RECT 20.5000 1370.5150 99.2650 1371.0850 ;
      RECT 900.5000 1369.2850 999.5000 1370.5150 ;
      RECT 20.5000 1369.2850 119.5000 1370.5150 ;
      RECT 920.5700 1368.7150 999.5000 1369.2850 ;
      RECT 900.5000 1368.7150 920.0000 1369.2850 ;
      RECT 99.8350 1368.7150 119.5000 1369.2850 ;
      RECT 20.5000 1368.7150 99.2650 1369.2850 ;
      RECT 900.5000 1367.4850 999.5000 1368.7150 ;
      RECT 20.5000 1367.4850 119.5000 1368.7150 ;
      RECT 920.5700 1366.9150 999.5000 1367.4850 ;
      RECT 900.5000 1366.9150 920.0000 1367.4850 ;
      RECT 99.8350 1366.9150 119.5000 1367.4850 ;
      RECT 20.5000 1366.9150 99.2650 1367.4850 ;
      RECT 900.5000 1365.6850 999.5000 1366.9150 ;
      RECT 20.5000 1365.6850 119.5000 1366.9150 ;
      RECT 920.5700 1365.1150 999.5000 1365.6850 ;
      RECT 900.5000 1365.1150 920.0000 1365.6850 ;
      RECT 99.8350 1365.1150 119.5000 1365.6850 ;
      RECT 20.5000 1365.1150 99.2650 1365.6850 ;
      RECT 900.5000 1363.8850 999.5000 1365.1150 ;
      RECT 20.5000 1363.8850 119.5000 1365.1150 ;
      RECT 920.5700 1363.3150 999.5000 1363.8850 ;
      RECT 900.5000 1363.3150 920.0000 1363.8850 ;
      RECT 99.8350 1363.3150 119.5000 1363.8850 ;
      RECT 20.5000 1363.3150 99.2650 1363.8850 ;
      RECT 900.5000 1362.0850 999.5000 1363.3150 ;
      RECT 20.5000 1362.0850 119.5000 1363.3150 ;
      RECT 920.5700 1361.5150 999.5000 1362.0850 ;
      RECT 900.5000 1361.5150 920.0000 1362.0850 ;
      RECT 99.8350 1361.5150 119.5000 1362.0850 ;
      RECT 20.5000 1361.5150 99.2650 1362.0850 ;
      RECT 900.5000 1360.2850 999.5000 1361.5150 ;
      RECT 20.5000 1360.2850 119.5000 1361.5150 ;
      RECT 920.5700 1359.7150 999.5000 1360.2850 ;
      RECT 900.5000 1359.7150 920.0000 1360.2850 ;
      RECT 99.8350 1359.7150 119.5000 1360.2850 ;
      RECT 20.5000 1359.7150 99.2650 1360.2850 ;
      RECT 900.5000 1358.4850 999.5000 1359.7150 ;
      RECT 20.5000 1358.4850 119.5000 1359.7150 ;
      RECT 920.5700 1357.9150 999.5000 1358.4850 ;
      RECT 900.5000 1357.9150 920.0000 1358.4850 ;
      RECT 99.8350 1357.9150 119.5000 1358.4850 ;
      RECT 20.5000 1357.9150 99.2650 1358.4850 ;
      RECT 900.5000 1356.6850 999.5000 1357.9150 ;
      RECT 20.5000 1356.6850 119.5000 1357.9150 ;
      RECT 920.5700 1356.1150 999.5000 1356.6850 ;
      RECT 900.5000 1356.1150 920.0000 1356.6850 ;
      RECT 99.8350 1356.1150 119.5000 1356.6850 ;
      RECT 20.5000 1356.1150 99.2650 1356.6850 ;
      RECT 900.5000 1354.8850 999.5000 1356.1150 ;
      RECT 20.5000 1354.8850 119.5000 1356.1150 ;
      RECT 920.5700 1354.3150 999.5000 1354.8850 ;
      RECT 900.5000 1354.3150 920.0000 1354.8850 ;
      RECT 99.8350 1354.3150 119.5000 1354.8850 ;
      RECT 20.5000 1354.3150 99.2650 1354.8850 ;
      RECT 900.5000 1353.0850 999.5000 1354.3150 ;
      RECT 20.5000 1353.0850 119.5000 1354.3150 ;
      RECT 920.5700 1352.5150 999.5000 1353.0850 ;
      RECT 900.5000 1352.5150 920.0000 1353.0850 ;
      RECT 99.8350 1352.5150 119.5000 1353.0850 ;
      RECT 20.5000 1352.5150 99.2650 1353.0850 ;
      RECT 900.5000 1351.2850 999.5000 1352.5150 ;
      RECT 20.5000 1351.2850 119.5000 1352.5150 ;
      RECT 920.5700 1350.7150 999.5000 1351.2850 ;
      RECT 900.5000 1350.7150 920.0000 1351.2850 ;
      RECT 99.8350 1350.7150 119.5000 1351.2850 ;
      RECT 20.5000 1350.7150 99.2650 1351.2850 ;
      RECT 900.5000 1349.4850 999.5000 1350.7150 ;
      RECT 20.5000 1349.4850 119.5000 1350.7150 ;
      RECT 920.5700 1348.9150 999.5000 1349.4850 ;
      RECT 900.5000 1348.9150 920.0000 1349.4850 ;
      RECT 99.8350 1348.9150 119.5000 1349.4850 ;
      RECT 20.5000 1348.9150 99.2650 1349.4850 ;
      RECT 900.5000 1347.6850 999.5000 1348.9150 ;
      RECT 20.5000 1347.6850 119.5000 1348.9150 ;
      RECT 920.5700 1347.1150 999.5000 1347.6850 ;
      RECT 900.5000 1347.1150 920.0000 1347.6850 ;
      RECT 99.8350 1347.1150 119.5000 1347.6850 ;
      RECT 20.5000 1347.1150 99.2650 1347.6850 ;
      RECT 900.5000 1345.8850 999.5000 1347.1150 ;
      RECT 20.5000 1345.8850 119.5000 1347.1150 ;
      RECT 920.5700 1345.3150 999.5000 1345.8850 ;
      RECT 900.5000 1345.3150 920.0000 1345.8850 ;
      RECT 99.8350 1345.3150 119.5000 1345.8850 ;
      RECT 20.5000 1345.3150 99.2650 1345.8850 ;
      RECT 900.5000 1344.0850 999.5000 1345.3150 ;
      RECT 20.5000 1344.0850 119.5000 1345.3150 ;
      RECT 920.5700 1343.5150 999.5000 1344.0850 ;
      RECT 900.5000 1343.5150 920.0000 1344.0850 ;
      RECT 99.8350 1343.5150 119.5000 1344.0850 ;
      RECT 20.5000 1343.5150 99.2650 1344.0850 ;
      RECT 900.5000 1342.2850 999.5000 1343.5150 ;
      RECT 20.5000 1342.2850 119.5000 1343.5150 ;
      RECT 920.5700 1341.7150 999.5000 1342.2850 ;
      RECT 900.5000 1341.7150 920.0000 1342.2850 ;
      RECT 99.8350 1341.7150 119.5000 1342.2850 ;
      RECT 20.5000 1341.7150 99.2650 1342.2850 ;
      RECT 900.5000 1340.4850 999.5000 1341.7150 ;
      RECT 20.5000 1340.4850 119.5000 1341.7150 ;
      RECT 920.5700 1339.9150 999.5000 1340.4850 ;
      RECT 900.5000 1339.9150 920.0000 1340.4850 ;
      RECT 99.8350 1339.9150 119.5000 1340.4850 ;
      RECT 20.5000 1339.9150 99.2650 1340.4850 ;
      RECT 900.5000 1338.6850 999.5000 1339.9150 ;
      RECT 20.5000 1338.6850 119.5000 1339.9150 ;
      RECT 920.5700 1338.1150 999.5000 1338.6850 ;
      RECT 900.5000 1338.1150 920.0000 1338.6850 ;
      RECT 99.8350 1338.1150 119.5000 1338.6850 ;
      RECT 20.5000 1338.1150 99.2650 1338.6850 ;
      RECT 900.5000 1336.8850 999.5000 1338.1150 ;
      RECT 20.5000 1336.8850 119.5000 1338.1150 ;
      RECT 920.5700 1336.3150 999.5000 1336.8850 ;
      RECT 900.5000 1336.3150 920.0000 1336.8850 ;
      RECT 99.8350 1336.3150 119.5000 1336.8850 ;
      RECT 20.5000 1336.3150 99.2650 1336.8850 ;
      RECT 900.5000 1335.0850 999.5000 1336.3150 ;
      RECT 20.5000 1335.0850 119.5000 1336.3150 ;
      RECT 920.5700 1334.5150 999.5000 1335.0850 ;
      RECT 900.5000 1334.5150 920.0000 1335.0850 ;
      RECT 99.8350 1334.5150 119.5000 1335.0850 ;
      RECT 20.5000 1334.5150 99.2650 1335.0850 ;
      RECT 900.5000 1333.2850 999.5000 1334.5150 ;
      RECT 20.5000 1333.2850 119.5000 1334.5150 ;
      RECT 920.5700 1332.7150 999.5000 1333.2850 ;
      RECT 900.5000 1332.7150 920.0000 1333.2850 ;
      RECT 99.8350 1332.7150 119.5000 1333.2850 ;
      RECT 20.5000 1332.7150 99.2650 1333.2850 ;
      RECT 900.5000 1331.4850 999.5000 1332.7150 ;
      RECT 20.5000 1331.4850 119.5000 1332.7150 ;
      RECT 920.5700 1330.9150 999.5000 1331.4850 ;
      RECT 900.5000 1330.9150 920.0000 1331.4850 ;
      RECT 99.8350 1330.9150 119.5000 1331.4850 ;
      RECT 20.5000 1330.9150 99.2650 1331.4850 ;
      RECT 900.5000 1329.6850 999.5000 1330.9150 ;
      RECT 20.5000 1329.6850 119.5000 1330.9150 ;
      RECT 920.5700 1329.1150 999.5000 1329.6850 ;
      RECT 900.5000 1329.1150 920.0000 1329.6850 ;
      RECT 99.8350 1329.1150 119.5000 1329.6850 ;
      RECT 20.5000 1329.1150 99.2650 1329.6850 ;
      RECT 900.5000 1327.8850 999.5000 1329.1150 ;
      RECT 20.5000 1327.8850 119.5000 1329.1150 ;
      RECT 920.5700 1327.3150 999.5000 1327.8850 ;
      RECT 900.5000 1327.3150 920.0000 1327.8850 ;
      RECT 99.8350 1327.3150 119.5000 1327.8850 ;
      RECT 20.5000 1327.3150 99.2650 1327.8850 ;
      RECT 900.5000 1326.0850 999.5000 1327.3150 ;
      RECT 20.5000 1326.0850 119.5000 1327.3150 ;
      RECT 920.5700 1325.5150 999.5000 1326.0850 ;
      RECT 900.5000 1325.5150 920.0000 1326.0850 ;
      RECT 99.8350 1325.5150 119.5000 1326.0850 ;
      RECT 20.5000 1325.5150 99.2650 1326.0850 ;
      RECT 900.5000 1324.2850 999.5000 1325.5150 ;
      RECT 20.5000 1324.2850 119.5000 1325.5150 ;
      RECT 920.5700 1323.7150 999.5000 1324.2850 ;
      RECT 900.5000 1323.7150 920.0000 1324.2850 ;
      RECT 99.8350 1323.7150 119.5000 1324.2850 ;
      RECT 20.5000 1323.7150 99.2650 1324.2850 ;
      RECT 900.5000 1322.4850 999.5000 1323.7150 ;
      RECT 20.5000 1322.4850 119.5000 1323.7150 ;
      RECT 920.5700 1321.9150 999.5000 1322.4850 ;
      RECT 900.5000 1321.9150 920.0000 1322.4850 ;
      RECT 99.8350 1321.9150 119.5000 1322.4850 ;
      RECT 20.5000 1321.9150 99.2650 1322.4850 ;
      RECT 900.5000 1320.6850 999.5000 1321.9150 ;
      RECT 20.5000 1320.6850 119.5000 1321.9150 ;
      RECT 920.5700 1320.1150 999.5000 1320.6850 ;
      RECT 900.5000 1320.1150 920.0000 1320.6850 ;
      RECT 99.8350 1320.1150 119.5000 1320.6850 ;
      RECT 20.5000 1320.1150 99.2650 1320.6850 ;
      RECT 900.5000 1318.8850 999.5000 1320.1150 ;
      RECT 20.5000 1318.8850 119.5000 1320.1150 ;
      RECT 920.5700 1318.3150 999.5000 1318.8850 ;
      RECT 900.5000 1318.3150 920.0000 1318.8850 ;
      RECT 99.8350 1318.3150 119.5000 1318.8850 ;
      RECT 20.5000 1318.3150 99.2650 1318.8850 ;
      RECT 900.5000 1317.0850 999.5000 1318.3150 ;
      RECT 20.5000 1317.0850 119.5000 1318.3150 ;
      RECT 920.5700 1316.5150 999.5000 1317.0850 ;
      RECT 900.5000 1316.5150 920.0000 1317.0850 ;
      RECT 99.8350 1316.5150 119.5000 1317.0850 ;
      RECT 20.5000 1316.5150 99.2650 1317.0850 ;
      RECT 900.5000 1315.2850 999.5000 1316.5150 ;
      RECT 20.5000 1315.2850 119.5000 1316.5150 ;
      RECT 920.5700 1314.7150 999.5000 1315.2850 ;
      RECT 900.5000 1314.7150 920.0000 1315.2850 ;
      RECT 99.8350 1314.7150 119.5000 1315.2850 ;
      RECT 20.5000 1314.7150 99.2650 1315.2850 ;
      RECT 900.5000 1313.4850 999.5000 1314.7150 ;
      RECT 20.5000 1313.4850 119.5000 1314.7150 ;
      RECT 920.5700 1312.9150 999.5000 1313.4850 ;
      RECT 900.5000 1312.9150 920.0000 1313.4850 ;
      RECT 99.8350 1312.9150 119.5000 1313.4850 ;
      RECT 20.5000 1312.9150 99.2650 1313.4850 ;
      RECT 900.5000 1311.6850 999.5000 1312.9150 ;
      RECT 20.5000 1311.6850 119.5000 1312.9150 ;
      RECT 920.5700 1311.1150 999.5000 1311.6850 ;
      RECT 900.5000 1311.1150 920.0000 1311.6850 ;
      RECT 99.8350 1311.1150 119.5000 1311.6850 ;
      RECT 20.5000 1311.1150 99.2650 1311.6850 ;
      RECT 900.5000 1309.8850 999.5000 1311.1150 ;
      RECT 20.5000 1309.8850 119.5000 1311.1150 ;
      RECT 920.5700 1309.3150 999.5000 1309.8850 ;
      RECT 900.5000 1309.3150 920.0000 1309.8850 ;
      RECT 99.8350 1309.3150 119.5000 1309.8850 ;
      RECT 20.5000 1309.3150 99.2650 1309.8850 ;
      RECT 900.5000 1308.0850 999.5000 1309.3150 ;
      RECT 20.5000 1308.0850 119.5000 1309.3150 ;
      RECT 920.5700 1307.5150 999.5000 1308.0850 ;
      RECT 900.5000 1307.5150 920.0000 1308.0850 ;
      RECT 99.8350 1307.5150 119.5000 1308.0850 ;
      RECT 20.5000 1307.5150 99.2650 1308.0850 ;
      RECT 900.5000 1306.2850 999.5000 1307.5150 ;
      RECT 20.5000 1306.2850 119.5000 1307.5150 ;
      RECT 920.5700 1305.7150 999.5000 1306.2850 ;
      RECT 900.5000 1305.7150 920.0000 1306.2850 ;
      RECT 99.8350 1305.7150 119.5000 1306.2850 ;
      RECT 20.5000 1305.7150 99.2650 1306.2850 ;
      RECT 900.5000 1304.4850 999.5000 1305.7150 ;
      RECT 20.5000 1304.4850 119.5000 1305.7150 ;
      RECT 920.5700 1303.9150 999.5000 1304.4850 ;
      RECT 900.5000 1303.9150 920.0000 1304.4850 ;
      RECT 99.8350 1303.9150 119.5000 1304.4850 ;
      RECT 20.5000 1303.9150 99.2650 1304.4850 ;
      RECT 900.5000 1302.6850 999.5000 1303.9150 ;
      RECT 20.5000 1302.6850 119.5000 1303.9150 ;
      RECT 920.5700 1302.1150 999.5000 1302.6850 ;
      RECT 900.5000 1302.1150 920.0000 1302.6850 ;
      RECT 99.8350 1302.1150 119.5000 1302.6850 ;
      RECT 20.5000 1302.1150 99.2650 1302.6850 ;
      RECT 900.5000 1300.8850 999.5000 1302.1150 ;
      RECT 20.5000 1300.8850 119.5000 1302.1150 ;
      RECT 920.5700 1300.3150 999.5000 1300.8850 ;
      RECT 900.5000 1300.3150 920.0000 1300.8850 ;
      RECT 99.8350 1300.3150 119.5000 1300.8850 ;
      RECT 20.5000 1300.3150 99.2650 1300.8850 ;
      RECT 900.5000 1299.0850 999.5000 1300.3150 ;
      RECT 20.5000 1299.0850 119.5000 1300.3150 ;
      RECT 920.5700 1298.5150 999.5000 1299.0850 ;
      RECT 900.5000 1298.5150 920.0000 1299.0850 ;
      RECT 99.8350 1298.5150 119.5000 1299.0850 ;
      RECT 20.5000 1298.5150 99.2650 1299.0850 ;
      RECT 900.5000 1297.2850 999.5000 1298.5150 ;
      RECT 20.5000 1297.2850 119.5000 1298.5150 ;
      RECT 920.5700 1296.7150 999.5000 1297.2850 ;
      RECT 900.5000 1296.7150 920.0000 1297.2850 ;
      RECT 99.8350 1296.7150 119.5000 1297.2850 ;
      RECT 20.5000 1296.7150 99.2650 1297.2850 ;
      RECT 900.5000 1295.4850 999.5000 1296.7150 ;
      RECT 20.5000 1295.4850 119.5000 1296.7150 ;
      RECT 920.5700 1294.9150 999.5000 1295.4850 ;
      RECT 900.5000 1294.9150 920.0000 1295.4850 ;
      RECT 99.8350 1294.9150 119.5000 1295.4850 ;
      RECT 20.5000 1294.9150 99.2650 1295.4850 ;
      RECT 900.5000 1293.6850 999.5000 1294.9150 ;
      RECT 20.5000 1293.6850 119.5000 1294.9150 ;
      RECT 920.5700 1293.1150 999.5000 1293.6850 ;
      RECT 900.5000 1293.1150 920.0000 1293.6850 ;
      RECT 99.8350 1293.1150 119.5000 1293.6850 ;
      RECT 20.5000 1293.1150 99.2650 1293.6850 ;
      RECT 900.5000 1291.8850 999.5000 1293.1150 ;
      RECT 20.5000 1291.8850 119.5000 1293.1150 ;
      RECT 920.5700 1291.3150 999.5000 1291.8850 ;
      RECT 900.5000 1291.3150 920.0000 1291.8850 ;
      RECT 99.8350 1291.3150 119.5000 1291.8850 ;
      RECT 20.5000 1291.3150 99.2650 1291.8850 ;
      RECT 900.5000 1290.0850 999.5000 1291.3150 ;
      RECT 20.5000 1290.0850 119.5000 1291.3150 ;
      RECT 920.5700 1289.5150 999.5000 1290.0850 ;
      RECT 900.5000 1289.5150 920.0000 1290.0850 ;
      RECT 99.8350 1289.5150 119.5000 1290.0850 ;
      RECT 20.5000 1289.5150 99.2650 1290.0850 ;
      RECT 900.5000 1288.2850 999.5000 1289.5150 ;
      RECT 20.5000 1288.2850 119.5000 1289.5150 ;
      RECT 920.5700 1287.7150 999.5000 1288.2850 ;
      RECT 900.5000 1287.7150 920.0000 1288.2850 ;
      RECT 99.8350 1287.7150 119.5000 1288.2850 ;
      RECT 20.5000 1287.7150 99.2650 1288.2850 ;
      RECT 900.5000 1286.4850 999.5000 1287.7150 ;
      RECT 20.5000 1286.4850 119.5000 1287.7150 ;
      RECT 920.5700 1285.9150 999.5000 1286.4850 ;
      RECT 900.5000 1285.9150 920.0000 1286.4850 ;
      RECT 99.8350 1285.9150 119.5000 1286.4850 ;
      RECT 20.5000 1285.9150 99.2650 1286.4850 ;
      RECT 900.5000 1284.6850 999.5000 1285.9150 ;
      RECT 20.5000 1284.6850 119.5000 1285.9150 ;
      RECT 920.5700 1284.1150 999.5000 1284.6850 ;
      RECT 900.5000 1284.1150 920.0000 1284.6850 ;
      RECT 99.8350 1284.1150 119.5000 1284.6850 ;
      RECT 20.5000 1284.1150 99.2650 1284.6850 ;
      RECT 900.5000 1282.8850 999.5000 1284.1150 ;
      RECT 20.5000 1282.8850 119.5000 1284.1150 ;
      RECT 920.5700 1282.3150 999.5000 1282.8850 ;
      RECT 900.5000 1282.3150 920.0000 1282.8850 ;
      RECT 99.8350 1282.3150 119.5000 1282.8850 ;
      RECT 20.5000 1282.3150 99.2650 1282.8850 ;
      RECT 900.5000 1281.0850 999.5000 1282.3150 ;
      RECT 20.5000 1281.0850 119.5000 1282.3150 ;
      RECT 920.5700 1280.5150 999.5000 1281.0850 ;
      RECT 900.5000 1280.5150 920.0000 1281.0850 ;
      RECT 99.8350 1280.5150 119.5000 1281.0850 ;
      RECT 20.5000 1280.5150 99.2650 1281.0850 ;
      RECT 900.5000 1279.2850 999.5000 1280.5150 ;
      RECT 20.5000 1279.2850 119.5000 1280.5150 ;
      RECT 920.5700 1278.7150 999.5000 1279.2850 ;
      RECT 900.5000 1278.7150 920.0000 1279.2850 ;
      RECT 99.8350 1278.7150 119.5000 1279.2850 ;
      RECT 20.5000 1278.7150 99.2650 1279.2850 ;
      RECT 900.5000 1277.4850 999.5000 1278.7150 ;
      RECT 20.5000 1277.4850 119.5000 1278.7150 ;
      RECT 920.5700 1276.9150 999.5000 1277.4850 ;
      RECT 900.5000 1276.9150 920.0000 1277.4850 ;
      RECT 99.8350 1276.9150 119.5000 1277.4850 ;
      RECT 20.5000 1276.9150 99.2650 1277.4850 ;
      RECT 900.5000 1275.6850 999.5000 1276.9150 ;
      RECT 20.5000 1275.6850 119.5000 1276.9150 ;
      RECT 920.5700 1275.1150 999.5000 1275.6850 ;
      RECT 900.5000 1275.1150 920.0000 1275.6850 ;
      RECT 99.8350 1275.1150 119.5000 1275.6850 ;
      RECT 20.5000 1275.1150 99.2650 1275.6850 ;
      RECT 900.5000 1273.8850 999.5000 1275.1150 ;
      RECT 20.5000 1273.8850 119.5000 1275.1150 ;
      RECT 920.5700 1273.3150 999.5000 1273.8850 ;
      RECT 900.5000 1273.3150 920.0000 1273.8850 ;
      RECT 99.8350 1273.3150 119.5000 1273.8850 ;
      RECT 20.5000 1273.3150 99.2650 1273.8850 ;
      RECT 900.5000 1272.0850 999.5000 1273.3150 ;
      RECT 20.5000 1272.0850 119.5000 1273.3150 ;
      RECT 920.5700 1271.5150 999.5000 1272.0850 ;
      RECT 900.5000 1271.5150 920.0000 1272.0850 ;
      RECT 99.8350 1271.5150 119.5000 1272.0850 ;
      RECT 20.5000 1271.5150 99.2650 1272.0850 ;
      RECT 900.5000 1270.2850 999.5000 1271.5150 ;
      RECT 20.5000 1270.2850 119.5000 1271.5150 ;
      RECT 920.5700 1269.7150 999.5000 1270.2850 ;
      RECT 900.5000 1269.7150 920.0000 1270.2850 ;
      RECT 99.8350 1269.7150 119.5000 1270.2850 ;
      RECT 20.5000 1269.7150 99.2650 1270.2850 ;
      RECT 900.5000 1268.4850 999.5000 1269.7150 ;
      RECT 20.5000 1268.4850 119.5000 1269.7150 ;
      RECT 920.5700 1267.9150 999.5000 1268.4850 ;
      RECT 900.5000 1267.9150 920.0000 1268.4850 ;
      RECT 99.8350 1267.9150 119.5000 1268.4850 ;
      RECT 20.5000 1267.9150 99.2650 1268.4850 ;
      RECT 900.5000 1266.6850 999.5000 1267.9150 ;
      RECT 20.5000 1266.6850 119.5000 1267.9150 ;
      RECT 920.5700 1266.1150 999.5000 1266.6850 ;
      RECT 900.5000 1266.1150 920.0000 1266.6850 ;
      RECT 99.8350 1266.1150 119.5000 1266.6850 ;
      RECT 20.5000 1266.1150 99.2650 1266.6850 ;
      RECT 900.5000 1264.8850 999.5000 1266.1150 ;
      RECT 20.5000 1264.8850 119.5000 1266.1150 ;
      RECT 920.5700 1264.3150 999.5000 1264.8850 ;
      RECT 900.5000 1264.3150 920.0000 1264.8850 ;
      RECT 99.8350 1264.3150 119.5000 1264.8850 ;
      RECT 20.5000 1264.3150 99.2650 1264.8850 ;
      RECT 900.5000 1263.0850 999.5000 1264.3150 ;
      RECT 20.5000 1263.0850 119.5000 1264.3150 ;
      RECT 920.5700 1262.5150 999.5000 1263.0850 ;
      RECT 900.5000 1262.5150 920.0000 1263.0850 ;
      RECT 99.8350 1262.5150 119.5000 1263.0850 ;
      RECT 20.5000 1262.5150 99.2650 1263.0850 ;
      RECT 900.5000 1261.2850 999.5000 1262.5150 ;
      RECT 20.5000 1261.2850 119.5000 1262.5150 ;
      RECT 920.5700 1260.7150 999.5000 1261.2850 ;
      RECT 900.5000 1260.7150 920.0000 1261.2850 ;
      RECT 99.8350 1260.7150 119.5000 1261.2850 ;
      RECT 20.5000 1260.7150 99.2650 1261.2850 ;
      RECT 900.5000 1259.4850 999.5000 1260.7150 ;
      RECT 20.5000 1259.4850 119.5000 1260.7150 ;
      RECT 920.5700 1258.9150 999.5000 1259.4850 ;
      RECT 900.5000 1258.9150 920.0000 1259.4850 ;
      RECT 99.8350 1258.9150 119.5000 1259.4850 ;
      RECT 20.5000 1258.9150 99.2650 1259.4850 ;
      RECT 900.5000 1257.6850 999.5000 1258.9150 ;
      RECT 20.5000 1257.6850 119.5000 1258.9150 ;
      RECT 920.5700 1257.1150 999.5000 1257.6850 ;
      RECT 900.5000 1257.1150 920.0000 1257.6850 ;
      RECT 99.8350 1257.1150 119.5000 1257.6850 ;
      RECT 20.5000 1257.1150 99.2650 1257.6850 ;
      RECT 900.5000 1255.8850 999.5000 1257.1150 ;
      RECT 20.5000 1255.8850 119.5000 1257.1150 ;
      RECT 920.5700 1255.3150 999.5000 1255.8850 ;
      RECT 900.5000 1255.3150 920.0000 1255.8850 ;
      RECT 99.8350 1255.3150 119.5000 1255.8850 ;
      RECT 20.5000 1255.3150 99.2650 1255.8850 ;
      RECT 900.5000 1254.0850 999.5000 1255.3150 ;
      RECT 20.5000 1254.0850 119.5000 1255.3150 ;
      RECT 920.5700 1253.5150 999.5000 1254.0850 ;
      RECT 900.5000 1253.5150 920.0000 1254.0850 ;
      RECT 99.8350 1253.5150 119.5000 1254.0850 ;
      RECT 20.5000 1253.5150 99.2650 1254.0850 ;
      RECT 900.5000 1252.2850 999.5000 1253.5150 ;
      RECT 20.5000 1252.2850 119.5000 1253.5150 ;
      RECT 920.5700 1251.7150 999.5000 1252.2850 ;
      RECT 900.5000 1251.7150 920.0000 1252.2850 ;
      RECT 99.8350 1251.7150 119.5000 1252.2850 ;
      RECT 20.5000 1251.7150 99.2650 1252.2850 ;
      RECT 900.5000 1250.4850 999.5000 1251.7150 ;
      RECT 20.5000 1250.4850 119.5000 1251.7150 ;
      RECT 920.5700 1249.9150 999.5000 1250.4850 ;
      RECT 900.5000 1249.9150 920.0000 1250.4850 ;
      RECT 99.8350 1249.9150 119.5000 1250.4850 ;
      RECT 20.5000 1249.9150 99.2650 1250.4850 ;
      RECT 900.5000 1248.6850 999.5000 1249.9150 ;
      RECT 20.5000 1248.6850 119.5000 1249.9150 ;
      RECT 920.5700 1248.1150 999.5000 1248.6850 ;
      RECT 900.5000 1248.1150 920.0000 1248.6850 ;
      RECT 99.8350 1248.1150 119.5000 1248.6850 ;
      RECT 20.5000 1248.1150 99.2650 1248.6850 ;
      RECT 900.5000 1246.8850 999.5000 1248.1150 ;
      RECT 20.5000 1246.8850 119.5000 1248.1150 ;
      RECT 920.5700 1246.3150 999.5000 1246.8850 ;
      RECT 900.5000 1246.3150 920.0000 1246.8850 ;
      RECT 99.8350 1246.3150 119.5000 1246.8850 ;
      RECT 20.5000 1246.3150 99.2650 1246.8850 ;
      RECT 900.5000 1245.0850 999.5000 1246.3150 ;
      RECT 20.5000 1245.0850 119.5000 1246.3150 ;
      RECT 920.5700 1244.5150 999.5000 1245.0850 ;
      RECT 900.5000 1244.5150 920.0000 1245.0850 ;
      RECT 99.8350 1244.5150 119.5000 1245.0850 ;
      RECT 20.5000 1244.5150 99.2650 1245.0850 ;
      RECT 900.5000 1243.2850 999.5000 1244.5150 ;
      RECT 20.5000 1243.2850 119.5000 1244.5150 ;
      RECT 920.5700 1242.7150 999.5000 1243.2850 ;
      RECT 900.5000 1242.7150 920.0000 1243.2850 ;
      RECT 99.8350 1242.7150 119.5000 1243.2850 ;
      RECT 20.5000 1242.7150 99.2650 1243.2850 ;
      RECT 900.5000 1241.4850 999.5000 1242.7150 ;
      RECT 20.5000 1241.4850 119.5000 1242.7150 ;
      RECT 920.5700 1240.9150 999.5000 1241.4850 ;
      RECT 900.5000 1240.9150 920.0000 1241.4850 ;
      RECT 99.8350 1240.9150 119.5000 1241.4850 ;
      RECT 20.5000 1240.9150 99.2650 1241.4850 ;
      RECT 900.5000 1239.6850 999.5000 1240.9150 ;
      RECT 20.5000 1239.6850 119.5000 1240.9150 ;
      RECT 920.5700 1239.1150 999.5000 1239.6850 ;
      RECT 900.5000 1239.1150 920.0000 1239.6850 ;
      RECT 99.8350 1239.1150 119.5000 1239.6850 ;
      RECT 20.5000 1239.1150 99.2650 1239.6850 ;
      RECT 900.5000 1237.8850 999.5000 1239.1150 ;
      RECT 20.5000 1237.8850 119.5000 1239.1150 ;
      RECT 920.5700 1237.3150 999.5000 1237.8850 ;
      RECT 900.5000 1237.3150 920.0000 1237.8850 ;
      RECT 99.8350 1237.3150 119.5000 1237.8850 ;
      RECT 20.5000 1237.3150 99.2650 1237.8850 ;
      RECT 900.5000 1236.0850 999.5000 1237.3150 ;
      RECT 20.5000 1236.0850 119.5000 1237.3150 ;
      RECT 920.5700 1235.5150 999.5000 1236.0850 ;
      RECT 900.5000 1235.5150 920.0000 1236.0850 ;
      RECT 99.8350 1235.5150 119.5000 1236.0850 ;
      RECT 20.5000 1235.5150 99.2650 1236.0850 ;
      RECT 900.5000 1234.2850 999.5000 1235.5150 ;
      RECT 20.5000 1234.2850 119.5000 1235.5150 ;
      RECT 920.5700 1233.7150 999.5000 1234.2850 ;
      RECT 900.5000 1233.7150 920.0000 1234.2850 ;
      RECT 99.8350 1233.7150 119.5000 1234.2850 ;
      RECT 20.5000 1233.7150 99.2650 1234.2850 ;
      RECT 900.5000 1232.4850 999.5000 1233.7150 ;
      RECT 20.5000 1232.4850 119.5000 1233.7150 ;
      RECT 920.5700 1231.9150 999.5000 1232.4850 ;
      RECT 900.5000 1231.9150 920.0000 1232.4850 ;
      RECT 99.8350 1231.9150 119.5000 1232.4850 ;
      RECT 20.5000 1231.9150 99.2650 1232.4850 ;
      RECT 900.5000 1230.6850 999.5000 1231.9150 ;
      RECT 20.5000 1230.6850 119.5000 1231.9150 ;
      RECT 920.5700 1230.1150 999.5000 1230.6850 ;
      RECT 900.5000 1230.1150 920.0000 1230.6850 ;
      RECT 99.8350 1230.1150 119.5000 1230.6850 ;
      RECT 20.5000 1230.1150 99.2650 1230.6850 ;
      RECT 900.5000 1228.8850 999.5000 1230.1150 ;
      RECT 20.5000 1228.8850 119.5000 1230.1150 ;
      RECT 920.5700 1228.3150 999.5000 1228.8850 ;
      RECT 900.5000 1228.3150 920.0000 1228.8850 ;
      RECT 99.8350 1228.3150 119.5000 1228.8850 ;
      RECT 20.5000 1228.3150 99.2650 1228.8850 ;
      RECT 900.5000 1227.0850 999.5000 1228.3150 ;
      RECT 20.5000 1227.0850 119.5000 1228.3150 ;
      RECT 920.5700 1226.5150 999.5000 1227.0850 ;
      RECT 900.5000 1226.5150 920.0000 1227.0850 ;
      RECT 99.8350 1226.5150 119.5000 1227.0850 ;
      RECT 20.5000 1226.5150 99.2650 1227.0850 ;
      RECT 900.5000 1225.2850 999.5000 1226.5150 ;
      RECT 20.5000 1225.2850 119.5000 1226.5150 ;
      RECT 920.5700 1224.7150 999.5000 1225.2850 ;
      RECT 900.5000 1224.7150 920.0000 1225.2850 ;
      RECT 99.8350 1224.7150 119.5000 1225.2850 ;
      RECT 20.5000 1224.7150 99.2650 1225.2850 ;
      RECT 900.5000 1223.4850 999.5000 1224.7150 ;
      RECT 20.5000 1223.4850 119.5000 1224.7150 ;
      RECT 920.5700 1222.9150 999.5000 1223.4850 ;
      RECT 900.5000 1222.9150 920.0000 1223.4850 ;
      RECT 99.8350 1222.9150 119.5000 1223.4850 ;
      RECT 20.5000 1222.9150 99.2650 1223.4850 ;
      RECT 900.5000 1221.6850 999.5000 1222.9150 ;
      RECT 20.5000 1221.6850 119.5000 1222.9150 ;
      RECT 920.5700 1221.1150 999.5000 1221.6850 ;
      RECT 900.5000 1221.1150 920.0000 1221.6850 ;
      RECT 99.8350 1221.1150 119.5000 1221.6850 ;
      RECT 20.5000 1221.1150 99.2650 1221.6850 ;
      RECT 900.5000 1219.8850 999.5000 1221.1150 ;
      RECT 20.5000 1219.8850 119.5000 1221.1150 ;
      RECT 920.5700 1219.3150 999.5000 1219.8850 ;
      RECT 900.5000 1219.3150 920.0000 1219.8850 ;
      RECT 99.8350 1219.3150 119.5000 1219.8850 ;
      RECT 20.5000 1219.3150 99.2650 1219.8850 ;
      RECT 900.5000 1218.0850 999.5000 1219.3150 ;
      RECT 20.5000 1218.0850 119.5000 1219.3150 ;
      RECT 920.5700 1217.5150 999.5000 1218.0850 ;
      RECT 900.5000 1217.5150 920.0000 1218.0850 ;
      RECT 99.8350 1217.5150 119.5000 1218.0850 ;
      RECT 20.5000 1217.5150 99.2650 1218.0850 ;
      RECT 900.5000 1216.2850 999.5000 1217.5150 ;
      RECT 20.5000 1216.2850 119.5000 1217.5150 ;
      RECT 920.5700 1215.7150 999.5000 1216.2850 ;
      RECT 900.5000 1215.7150 920.0000 1216.2850 ;
      RECT 99.8350 1215.7150 119.5000 1216.2850 ;
      RECT 20.5000 1215.7150 99.2650 1216.2850 ;
      RECT 900.5000 1214.4850 999.5000 1215.7150 ;
      RECT 20.5000 1214.4850 119.5000 1215.7150 ;
      RECT 920.5700 1213.9150 999.5000 1214.4850 ;
      RECT 900.5000 1213.9150 920.0000 1214.4850 ;
      RECT 99.8350 1213.9150 119.5000 1214.4850 ;
      RECT 20.5000 1213.9150 99.2650 1214.4850 ;
      RECT 900.5000 1212.6850 999.5000 1213.9150 ;
      RECT 20.5000 1212.6850 119.5000 1213.9150 ;
      RECT 920.5700 1212.1150 999.5000 1212.6850 ;
      RECT 900.5000 1212.1150 920.0000 1212.6850 ;
      RECT 99.8350 1212.1150 119.5000 1212.6850 ;
      RECT 20.5000 1212.1150 99.2650 1212.6850 ;
      RECT 900.5000 1210.8850 999.5000 1212.1150 ;
      RECT 20.5000 1210.8850 119.5000 1212.1150 ;
      RECT 920.5700 1210.3150 999.5000 1210.8850 ;
      RECT 900.5000 1210.3150 920.0000 1210.8850 ;
      RECT 99.8350 1210.3150 119.5000 1210.8850 ;
      RECT 20.5000 1210.3150 99.2650 1210.8850 ;
      RECT 900.5000 1209.0850 999.5000 1210.3150 ;
      RECT 20.5000 1209.0850 119.5000 1210.3150 ;
      RECT 920.5700 1208.5150 999.5000 1209.0850 ;
      RECT 900.5000 1208.5150 920.0000 1209.0850 ;
      RECT 99.8350 1208.5150 119.5000 1209.0850 ;
      RECT 20.5000 1208.5150 99.2650 1209.0850 ;
      RECT 900.5000 1207.2850 999.5000 1208.5150 ;
      RECT 20.5000 1207.2850 119.5000 1208.5150 ;
      RECT 920.5700 1206.7150 999.5000 1207.2850 ;
      RECT 900.5000 1206.7150 920.0000 1207.2850 ;
      RECT 99.8350 1206.7150 119.5000 1207.2850 ;
      RECT 20.5000 1206.7150 99.2650 1207.2850 ;
      RECT 900.5000 1205.4850 999.5000 1206.7150 ;
      RECT 20.5000 1205.4850 119.5000 1206.7150 ;
      RECT 920.5700 1204.9150 999.5000 1205.4850 ;
      RECT 900.5000 1204.9150 920.0000 1205.4850 ;
      RECT 99.8350 1204.9150 119.5000 1205.4850 ;
      RECT 20.5000 1204.9150 99.2650 1205.4850 ;
      RECT 900.5000 1203.6850 999.5000 1204.9150 ;
      RECT 20.5000 1203.6850 119.5000 1204.9150 ;
      RECT 920.5700 1203.1150 999.5000 1203.6850 ;
      RECT 900.5000 1203.1150 920.0000 1203.6850 ;
      RECT 99.8350 1203.1150 119.5000 1203.6850 ;
      RECT 20.5000 1203.1150 99.2650 1203.6850 ;
      RECT 900.5000 1201.8850 999.5000 1203.1150 ;
      RECT 20.5000 1201.8850 119.5000 1203.1150 ;
      RECT 920.5700 1201.3150 999.5000 1201.8850 ;
      RECT 900.5000 1201.3150 920.0000 1201.8850 ;
      RECT 99.8350 1201.3150 119.5000 1201.8850 ;
      RECT 20.5000 1201.3150 99.2650 1201.8850 ;
      RECT 900.5000 1200.0850 999.5000 1201.3150 ;
      RECT 20.5000 1200.0850 119.5000 1201.3150 ;
      RECT 920.5700 1199.5150 999.5000 1200.0850 ;
      RECT 900.5000 1199.5150 920.0000 1200.0850 ;
      RECT 99.8350 1199.5150 119.5000 1200.0850 ;
      RECT 20.5000 1199.5150 99.2650 1200.0850 ;
      RECT 900.5000 1198.2850 999.5000 1199.5150 ;
      RECT 20.5000 1198.2850 119.5000 1199.5150 ;
      RECT 920.5700 1197.7150 999.5000 1198.2850 ;
      RECT 900.5000 1197.7150 920.0000 1198.2850 ;
      RECT 99.8350 1197.7150 119.5000 1198.2850 ;
      RECT 20.5000 1197.7150 99.2650 1198.2850 ;
      RECT 900.5000 1196.4850 999.5000 1197.7150 ;
      RECT 20.5000 1196.4850 119.5000 1197.7150 ;
      RECT 920.5700 1195.9150 999.5000 1196.4850 ;
      RECT 900.5000 1195.9150 920.0000 1196.4850 ;
      RECT 99.8350 1195.9150 119.5000 1196.4850 ;
      RECT 20.5000 1195.9150 99.2650 1196.4850 ;
      RECT 900.5000 1194.6850 999.5000 1195.9150 ;
      RECT 20.5000 1194.6850 119.5000 1195.9150 ;
      RECT 920.5700 1194.1150 999.5000 1194.6850 ;
      RECT 900.5000 1194.1150 920.0000 1194.6850 ;
      RECT 99.8350 1194.1150 119.5000 1194.6850 ;
      RECT 20.5000 1194.1150 99.2650 1194.6850 ;
      RECT 900.5000 1192.8850 999.5000 1194.1150 ;
      RECT 20.5000 1192.8850 119.5000 1194.1150 ;
      RECT 920.5700 1192.3150 999.5000 1192.8850 ;
      RECT 900.5000 1192.3150 920.0000 1192.8850 ;
      RECT 99.8350 1192.3150 119.5000 1192.8850 ;
      RECT 20.5000 1192.3150 99.2650 1192.8850 ;
      RECT 900.5000 1191.0850 999.5000 1192.3150 ;
      RECT 20.5000 1191.0850 119.5000 1192.3150 ;
      RECT 920.5700 1190.5150 999.5000 1191.0850 ;
      RECT 900.5000 1190.5150 920.0000 1191.0850 ;
      RECT 99.8350 1190.5150 119.5000 1191.0850 ;
      RECT 20.5000 1190.5150 99.2650 1191.0850 ;
      RECT 900.5000 1189.2850 999.5000 1190.5150 ;
      RECT 20.5000 1189.2850 119.5000 1190.5150 ;
      RECT 920.5700 1188.7150 999.5000 1189.2850 ;
      RECT 900.5000 1188.7150 920.0000 1189.2850 ;
      RECT 99.8350 1188.7150 119.5000 1189.2850 ;
      RECT 20.5000 1188.7150 99.2650 1189.2850 ;
      RECT 900.5000 1187.4850 999.5000 1188.7150 ;
      RECT 20.5000 1187.4850 119.5000 1188.7150 ;
      RECT 920.5700 1186.9150 999.5000 1187.4850 ;
      RECT 900.5000 1186.9150 920.0000 1187.4850 ;
      RECT 99.8350 1186.9150 119.5000 1187.4850 ;
      RECT 20.5000 1186.9150 99.2650 1187.4850 ;
      RECT 900.5000 1185.6850 999.5000 1186.9150 ;
      RECT 20.5000 1185.6850 119.5000 1186.9150 ;
      RECT 920.5700 1185.1150 999.5000 1185.6850 ;
      RECT 900.5000 1185.1150 920.0000 1185.6850 ;
      RECT 99.8350 1185.1150 119.5000 1185.6850 ;
      RECT 20.5000 1185.1150 99.2650 1185.6850 ;
      RECT 900.5000 1183.8850 999.5000 1185.1150 ;
      RECT 20.5000 1183.8850 119.5000 1185.1150 ;
      RECT 920.5700 1183.3150 999.5000 1183.8850 ;
      RECT 900.5000 1183.3150 920.0000 1183.8850 ;
      RECT 99.8350 1183.3150 119.5000 1183.8850 ;
      RECT 20.5000 1183.3150 99.2650 1183.8850 ;
      RECT 900.5000 1182.0850 999.5000 1183.3150 ;
      RECT 20.5000 1182.0850 119.5000 1183.3150 ;
      RECT 920.5700 1181.5150 999.5000 1182.0850 ;
      RECT 900.5000 1181.5150 920.0000 1182.0850 ;
      RECT 99.8350 1181.5150 119.5000 1182.0850 ;
      RECT 20.5000 1181.5150 99.2650 1182.0850 ;
      RECT 900.5000 1180.2850 999.5000 1181.5150 ;
      RECT 20.5000 1180.2850 119.5000 1181.5150 ;
      RECT 920.5700 1179.7150 999.5000 1180.2850 ;
      RECT 900.5000 1179.7150 920.0000 1180.2850 ;
      RECT 99.8350 1179.7150 119.5000 1180.2850 ;
      RECT 20.5000 1179.7150 99.2650 1180.2850 ;
      RECT 900.5000 1178.4850 999.5000 1179.7150 ;
      RECT 20.5000 1178.4850 119.5000 1179.7150 ;
      RECT 920.5700 1177.9150 999.5000 1178.4850 ;
      RECT 900.5000 1177.9150 920.0000 1178.4850 ;
      RECT 99.8350 1177.9150 119.5000 1178.4850 ;
      RECT 20.5000 1177.9150 99.2650 1178.4850 ;
      RECT 900.5000 1176.6850 999.5000 1177.9150 ;
      RECT 20.5000 1176.6850 119.5000 1177.9150 ;
      RECT 920.5700 1176.1150 999.5000 1176.6850 ;
      RECT 900.5000 1176.1150 920.0000 1176.6850 ;
      RECT 99.8350 1176.1150 119.5000 1176.6850 ;
      RECT 20.5000 1176.1150 99.2650 1176.6850 ;
      RECT 900.5000 1174.8850 999.5000 1176.1150 ;
      RECT 20.5000 1174.8850 119.5000 1176.1150 ;
      RECT 920.5700 1174.3150 999.5000 1174.8850 ;
      RECT 900.5000 1174.3150 920.0000 1174.8850 ;
      RECT 99.8350 1174.3150 119.5000 1174.8850 ;
      RECT 20.5000 1174.3150 99.2650 1174.8850 ;
      RECT 900.5000 1173.0850 999.5000 1174.3150 ;
      RECT 20.5000 1173.0850 119.5000 1174.3150 ;
      RECT 920.5700 1172.5150 999.5000 1173.0850 ;
      RECT 900.5000 1172.5150 920.0000 1173.0850 ;
      RECT 99.8350 1172.5150 119.5000 1173.0850 ;
      RECT 20.5000 1172.5150 99.2650 1173.0850 ;
      RECT 900.5000 1171.2850 999.5000 1172.5150 ;
      RECT 20.5000 1171.2850 119.5000 1172.5150 ;
      RECT 920.5700 1170.7150 999.5000 1171.2850 ;
      RECT 900.5000 1170.7150 920.0000 1171.2850 ;
      RECT 99.8350 1170.7150 119.5000 1171.2850 ;
      RECT 20.5000 1170.7150 99.2650 1171.2850 ;
      RECT 900.5000 1169.4850 999.5000 1170.7150 ;
      RECT 20.5000 1169.4850 119.5000 1170.7150 ;
      RECT 920.5700 1168.9150 999.5000 1169.4850 ;
      RECT 900.5000 1168.9150 920.0000 1169.4850 ;
      RECT 99.8350 1168.9150 119.5000 1169.4850 ;
      RECT 20.5000 1168.9150 99.2650 1169.4850 ;
      RECT 900.5000 1167.6850 999.5000 1168.9150 ;
      RECT 20.5000 1167.6850 119.5000 1168.9150 ;
      RECT 920.5700 1167.1150 999.5000 1167.6850 ;
      RECT 900.5000 1167.1150 920.0000 1167.6850 ;
      RECT 99.8350 1167.1150 119.5000 1167.6850 ;
      RECT 20.5000 1167.1150 99.2650 1167.6850 ;
      RECT 900.5000 1165.8850 999.5000 1167.1150 ;
      RECT 20.5000 1165.8850 119.5000 1167.1150 ;
      RECT 920.5700 1165.3150 999.5000 1165.8850 ;
      RECT 900.5000 1165.3150 920.0000 1165.8850 ;
      RECT 99.8350 1165.3150 119.5000 1165.8850 ;
      RECT 20.5000 1165.3150 99.2650 1165.8850 ;
      RECT 900.5000 1164.0850 999.5000 1165.3150 ;
      RECT 20.5000 1164.0850 119.5000 1165.3150 ;
      RECT 920.5700 1163.5150 999.5000 1164.0850 ;
      RECT 900.5000 1163.5150 920.0000 1164.0850 ;
      RECT 99.8350 1163.5150 119.5000 1164.0850 ;
      RECT 20.5000 1163.5150 99.2650 1164.0850 ;
      RECT 900.5000 1162.2850 999.5000 1163.5150 ;
      RECT 20.5000 1162.2850 119.5000 1163.5150 ;
      RECT 920.5700 1161.7150 999.5000 1162.2850 ;
      RECT 900.5000 1161.7150 920.0000 1162.2850 ;
      RECT 99.8350 1161.7150 119.5000 1162.2850 ;
      RECT 20.5000 1161.7150 99.2650 1162.2850 ;
      RECT 900.5000 1160.4850 999.5000 1161.7150 ;
      RECT 20.5000 1160.4850 119.5000 1161.7150 ;
      RECT 920.5700 1159.9150 999.5000 1160.4850 ;
      RECT 900.5000 1159.9150 920.0000 1160.4850 ;
      RECT 99.8350 1159.9150 119.5000 1160.4850 ;
      RECT 20.5000 1159.9150 99.2650 1160.4850 ;
      RECT 900.5000 1158.6850 999.5000 1159.9150 ;
      RECT 20.5000 1158.6850 119.5000 1159.9150 ;
      RECT 920.5700 1158.1150 999.5000 1158.6850 ;
      RECT 900.5000 1158.1150 920.0000 1158.6850 ;
      RECT 99.8350 1158.1150 119.5000 1158.6850 ;
      RECT 20.5000 1158.1150 99.2650 1158.6850 ;
      RECT 900.5000 1156.8850 999.5000 1158.1150 ;
      RECT 20.5000 1156.8850 119.5000 1158.1150 ;
      RECT 920.5700 1156.3150 999.5000 1156.8850 ;
      RECT 900.5000 1156.3150 920.0000 1156.8850 ;
      RECT 99.8350 1156.3150 119.5000 1156.8850 ;
      RECT 20.5000 1156.3150 99.2650 1156.8850 ;
      RECT 900.5000 1155.0850 999.5000 1156.3150 ;
      RECT 20.5000 1155.0850 119.5000 1156.3150 ;
      RECT 920.5700 1154.5150 999.5000 1155.0850 ;
      RECT 900.5000 1154.5150 920.0000 1155.0850 ;
      RECT 99.8350 1154.5150 119.5000 1155.0850 ;
      RECT 20.5000 1154.5150 99.2650 1155.0850 ;
      RECT 900.5000 1153.2850 999.5000 1154.5150 ;
      RECT 20.5000 1153.2850 119.5000 1154.5150 ;
      RECT 920.5700 1152.7150 999.5000 1153.2850 ;
      RECT 900.5000 1152.7150 920.0000 1153.2850 ;
      RECT 99.8350 1152.7150 119.5000 1153.2850 ;
      RECT 20.5000 1152.7150 99.2650 1153.2850 ;
      RECT 900.5000 1151.4850 999.5000 1152.7150 ;
      RECT 20.5000 1151.4850 119.5000 1152.7150 ;
      RECT 920.5700 1150.9150 999.5000 1151.4850 ;
      RECT 900.5000 1150.9150 920.0000 1151.4850 ;
      RECT 99.8350 1150.9150 119.5000 1151.4850 ;
      RECT 20.5000 1150.9150 99.2650 1151.4850 ;
      RECT 900.5000 1149.6850 999.5000 1150.9150 ;
      RECT 20.5000 1149.6850 119.5000 1150.9150 ;
      RECT 920.5700 1149.1150 999.5000 1149.6850 ;
      RECT 900.5000 1149.1150 920.0000 1149.6850 ;
      RECT 99.8350 1149.1150 119.5000 1149.6850 ;
      RECT 20.5000 1149.1150 99.2650 1149.6850 ;
      RECT 900.5000 1147.8850 999.5000 1149.1150 ;
      RECT 20.5000 1147.8850 119.5000 1149.1150 ;
      RECT 920.5700 1147.3150 999.5000 1147.8850 ;
      RECT 900.5000 1147.3150 920.0000 1147.8850 ;
      RECT 99.8350 1147.3150 119.5000 1147.8850 ;
      RECT 20.5000 1147.3150 99.2650 1147.8850 ;
      RECT 900.5000 1146.0850 999.5000 1147.3150 ;
      RECT 20.5000 1146.0850 119.5000 1147.3150 ;
      RECT 920.5700 1145.5150 999.5000 1146.0850 ;
      RECT 900.5000 1145.5150 920.0000 1146.0850 ;
      RECT 99.8350 1145.5150 119.5000 1146.0850 ;
      RECT 20.5000 1145.5150 99.2650 1146.0850 ;
      RECT 900.5000 1144.2850 999.5000 1145.5150 ;
      RECT 20.5000 1144.2850 119.5000 1145.5150 ;
      RECT 920.5700 1143.7150 999.5000 1144.2850 ;
      RECT 900.5000 1143.7150 920.0000 1144.2850 ;
      RECT 99.8350 1143.7150 119.5000 1144.2850 ;
      RECT 20.5000 1143.7150 99.2650 1144.2850 ;
      RECT 900.5000 1142.4850 999.5000 1143.7150 ;
      RECT 20.5000 1142.4850 119.5000 1143.7150 ;
      RECT 920.5700 1141.9150 999.5000 1142.4850 ;
      RECT 900.5000 1141.9150 920.0000 1142.4850 ;
      RECT 99.8350 1141.9150 119.5000 1142.4850 ;
      RECT 20.5000 1141.9150 99.2650 1142.4850 ;
      RECT 900.5000 1140.6850 999.5000 1141.9150 ;
      RECT 20.5000 1140.6850 119.5000 1141.9150 ;
      RECT 920.5700 1140.1150 999.5000 1140.6850 ;
      RECT 900.5000 1140.1150 920.0000 1140.6850 ;
      RECT 99.8350 1140.1150 119.5000 1140.6850 ;
      RECT 20.5000 1140.1150 99.2650 1140.6850 ;
      RECT 900.5000 1138.8850 999.5000 1140.1150 ;
      RECT 20.5000 1138.8850 119.5000 1140.1150 ;
      RECT 920.5700 1138.3150 999.5000 1138.8850 ;
      RECT 900.5000 1138.3150 920.0000 1138.8850 ;
      RECT 99.8350 1138.3150 119.5000 1138.8850 ;
      RECT 20.5000 1138.3150 99.2650 1138.8850 ;
      RECT 900.5000 1137.0850 999.5000 1138.3150 ;
      RECT 20.5000 1137.0850 119.5000 1138.3150 ;
      RECT 920.5700 1136.5150 999.5000 1137.0850 ;
      RECT 900.5000 1136.5150 920.0000 1137.0850 ;
      RECT 99.8350 1136.5150 119.5000 1137.0850 ;
      RECT 20.5000 1136.5150 99.2650 1137.0850 ;
      RECT 900.5000 1135.2850 999.5000 1136.5150 ;
      RECT 20.5000 1135.2850 119.5000 1136.5150 ;
      RECT 920.5700 1134.7150 999.5000 1135.2850 ;
      RECT 900.5000 1134.7150 920.0000 1135.2850 ;
      RECT 99.8350 1134.7150 119.5000 1135.2850 ;
      RECT 20.5000 1134.7150 99.2650 1135.2850 ;
      RECT 900.5000 1133.4850 999.5000 1134.7150 ;
      RECT 20.5000 1133.4850 119.5000 1134.7150 ;
      RECT 920.5700 1132.9150 999.5000 1133.4850 ;
      RECT 900.5000 1132.9150 920.0000 1133.4850 ;
      RECT 99.8350 1132.9150 119.5000 1133.4850 ;
      RECT 20.5000 1132.9150 99.2650 1133.4850 ;
      RECT 900.5000 1131.6850 999.5000 1132.9150 ;
      RECT 20.5000 1131.6850 119.5000 1132.9150 ;
      RECT 920.5700 1131.1150 999.5000 1131.6850 ;
      RECT 900.5000 1131.1150 920.0000 1131.6850 ;
      RECT 99.8350 1131.1150 119.5000 1131.6850 ;
      RECT 20.5000 1131.1150 99.2650 1131.6850 ;
      RECT 900.5000 1129.8850 999.5000 1131.1150 ;
      RECT 20.5000 1129.8850 119.5000 1131.1150 ;
      RECT 920.5700 1129.3150 999.5000 1129.8850 ;
      RECT 900.5000 1129.3150 920.0000 1129.8850 ;
      RECT 99.8350 1129.3150 119.5000 1129.8850 ;
      RECT 20.5000 1129.3150 99.2650 1129.8850 ;
      RECT 900.5000 1128.0850 999.5000 1129.3150 ;
      RECT 20.5000 1128.0850 119.5000 1129.3150 ;
      RECT 920.5700 1127.5150 999.5000 1128.0850 ;
      RECT 900.5000 1127.5150 920.0000 1128.0850 ;
      RECT 99.8350 1127.5150 119.5000 1128.0850 ;
      RECT 20.5000 1127.5150 99.2650 1128.0850 ;
      RECT 900.5000 1126.2850 999.5000 1127.5150 ;
      RECT 20.5000 1126.2850 119.5000 1127.5150 ;
      RECT 920.5700 1125.7150 999.5000 1126.2850 ;
      RECT 900.5000 1125.7150 920.0000 1126.2850 ;
      RECT 99.8350 1125.7150 119.5000 1126.2850 ;
      RECT 20.5000 1125.7150 99.2650 1126.2850 ;
      RECT 900.5000 1124.4850 999.5000 1125.7150 ;
      RECT 20.5000 1124.4850 119.5000 1125.7150 ;
      RECT 920.5700 1123.9150 999.5000 1124.4850 ;
      RECT 900.5000 1123.9150 920.0000 1124.4850 ;
      RECT 99.8350 1123.9150 119.5000 1124.4850 ;
      RECT 20.5000 1123.9150 99.2650 1124.4850 ;
      RECT 900.5000 1122.6850 999.5000 1123.9150 ;
      RECT 20.5000 1122.6850 119.5000 1123.9150 ;
      RECT 920.5700 1122.1150 999.5000 1122.6850 ;
      RECT 900.5000 1122.1150 920.0000 1122.6850 ;
      RECT 99.8350 1122.1150 119.5000 1122.6850 ;
      RECT 20.5000 1122.1150 99.2650 1122.6850 ;
      RECT 900.5000 1120.8850 999.5000 1122.1150 ;
      RECT 20.5000 1120.8850 119.5000 1122.1150 ;
      RECT 920.5700 1120.3150 999.5000 1120.8850 ;
      RECT 900.5000 1120.3150 920.0000 1120.8850 ;
      RECT 99.8350 1120.3150 119.5000 1120.8850 ;
      RECT 20.5000 1120.3150 99.2650 1120.8850 ;
      RECT 900.5000 1119.0850 999.5000 1120.3150 ;
      RECT 20.5000 1119.0850 119.5000 1120.3150 ;
      RECT 920.5700 1118.5150 999.5000 1119.0850 ;
      RECT 900.5000 1118.5150 920.0000 1119.0850 ;
      RECT 99.8350 1118.5150 119.5000 1119.0850 ;
      RECT 20.5000 1118.5150 99.2650 1119.0850 ;
      RECT 900.5000 1117.2850 999.5000 1118.5150 ;
      RECT 20.5000 1117.2850 119.5000 1118.5150 ;
      RECT 920.5700 1116.7150 999.5000 1117.2850 ;
      RECT 900.5000 1116.7150 920.0000 1117.2850 ;
      RECT 99.8350 1116.7150 119.5000 1117.2850 ;
      RECT 20.5000 1116.7150 99.2650 1117.2850 ;
      RECT 900.5000 1115.4850 999.5000 1116.7150 ;
      RECT 20.5000 1115.4850 119.5000 1116.7150 ;
      RECT 920.5700 1114.9150 999.5000 1115.4850 ;
      RECT 900.5000 1114.9150 920.0000 1115.4850 ;
      RECT 99.8350 1114.9150 119.5000 1115.4850 ;
      RECT 20.5000 1114.9150 99.2650 1115.4850 ;
      RECT 900.5000 1113.6850 999.5000 1114.9150 ;
      RECT 20.5000 1113.6850 119.5000 1114.9150 ;
      RECT 920.5700 1113.1150 999.5000 1113.6850 ;
      RECT 900.5000 1113.1150 920.0000 1113.6850 ;
      RECT 99.8350 1113.1150 119.5000 1113.6850 ;
      RECT 20.5000 1113.1150 99.2650 1113.6850 ;
      RECT 900.5000 1111.8850 999.5000 1113.1150 ;
      RECT 20.5000 1111.8850 119.5000 1113.1150 ;
      RECT 920.5700 1111.3150 999.5000 1111.8850 ;
      RECT 900.5000 1111.3150 920.0000 1111.8850 ;
      RECT 99.8350 1111.3150 119.5000 1111.8850 ;
      RECT 20.5000 1111.3150 99.2650 1111.8850 ;
      RECT 900.5000 1110.0850 999.5000 1111.3150 ;
      RECT 20.5000 1110.0850 119.5000 1111.3150 ;
      RECT 920.5700 1109.5150 999.5000 1110.0850 ;
      RECT 900.5000 1109.5150 920.0000 1110.0850 ;
      RECT 99.8350 1109.5150 119.5000 1110.0850 ;
      RECT 20.5000 1109.5150 99.2650 1110.0850 ;
      RECT 900.5000 1108.2850 999.5000 1109.5150 ;
      RECT 20.5000 1108.2850 119.5000 1109.5150 ;
      RECT 920.5700 1107.7150 999.5000 1108.2850 ;
      RECT 900.5000 1107.7150 920.0000 1108.2850 ;
      RECT 99.8350 1107.7150 119.5000 1108.2850 ;
      RECT 20.5000 1107.7150 99.2650 1108.2850 ;
      RECT 900.5000 1106.4850 999.5000 1107.7150 ;
      RECT 20.5000 1106.4850 119.5000 1107.7150 ;
      RECT 920.5700 1105.9150 999.5000 1106.4850 ;
      RECT 900.5000 1105.9150 920.0000 1106.4850 ;
      RECT 99.8350 1105.9150 119.5000 1106.4850 ;
      RECT 20.5000 1105.9150 99.2650 1106.4850 ;
      RECT 900.5000 1104.6850 999.5000 1105.9150 ;
      RECT 20.5000 1104.6850 119.5000 1105.9150 ;
      RECT 920.5700 1104.1150 999.5000 1104.6850 ;
      RECT 900.5000 1104.1150 920.0000 1104.6850 ;
      RECT 99.8350 1104.1150 119.5000 1104.6850 ;
      RECT 20.5000 1104.1150 99.2650 1104.6850 ;
      RECT 900.5000 1102.8850 999.5000 1104.1150 ;
      RECT 20.5000 1102.8850 119.5000 1104.1150 ;
      RECT 920.5700 1102.3150 999.5000 1102.8850 ;
      RECT 900.5000 1102.3150 920.0000 1102.8850 ;
      RECT 99.8350 1102.3150 119.5000 1102.8850 ;
      RECT 20.5000 1102.3150 99.2650 1102.8850 ;
      RECT 900.5000 1101.0850 999.5000 1102.3150 ;
      RECT 20.5000 1101.0850 119.5000 1102.3150 ;
      RECT 920.5700 1100.5150 999.5000 1101.0850 ;
      RECT 900.5000 1100.5150 920.0000 1101.0850 ;
      RECT 99.8350 1100.5150 119.5000 1101.0850 ;
      RECT 20.5000 1100.5150 99.2650 1101.0850 ;
      RECT 900.5000 1020.0850 999.5000 1100.5150 ;
      RECT 20.5000 1020.0850 119.5000 1100.5150 ;
      RECT 920.5700 1019.5150 999.5000 1020.0850 ;
      RECT 900.5000 1019.5150 920.0000 1020.0850 ;
      RECT 99.8350 1019.5150 119.5000 1020.0850 ;
      RECT 20.5000 1019.5150 99.2650 1020.0850 ;
      RECT 900.5000 1018.2850 999.5000 1019.5150 ;
      RECT 20.5000 1018.2850 119.5000 1019.5150 ;
      RECT 920.5700 1017.7150 999.5000 1018.2850 ;
      RECT 900.5000 1017.7150 920.0000 1018.2850 ;
      RECT 99.8350 1017.7150 119.5000 1018.2850 ;
      RECT 20.5000 1017.7150 99.2650 1018.2850 ;
      RECT 900.5000 1016.4850 999.5000 1017.7150 ;
      RECT 20.5000 1016.4850 119.5000 1017.7150 ;
      RECT 920.5700 1015.9150 999.5000 1016.4850 ;
      RECT 900.5000 1015.9150 920.0000 1016.4850 ;
      RECT 99.8350 1015.9150 119.5000 1016.4850 ;
      RECT 20.5000 1015.9150 99.2650 1016.4850 ;
      RECT 900.5000 1014.6850 999.5000 1015.9150 ;
      RECT 20.5000 1014.6850 119.5000 1015.9150 ;
      RECT 920.5700 1014.1150 999.5000 1014.6850 ;
      RECT 900.5000 1014.1150 920.0000 1014.6850 ;
      RECT 99.8350 1014.1150 119.5000 1014.6850 ;
      RECT 20.5000 1014.1150 99.2650 1014.6850 ;
      RECT 900.5000 1012.8850 999.5000 1014.1150 ;
      RECT 20.5000 1012.8850 119.5000 1014.1150 ;
      RECT 920.5700 1012.3150 999.5000 1012.8850 ;
      RECT 900.5000 1012.3150 920.0000 1012.8850 ;
      RECT 99.8350 1012.3150 119.5000 1012.8850 ;
      RECT 20.5000 1012.3150 99.2650 1012.8850 ;
      RECT 900.5000 1011.0850 999.5000 1012.3150 ;
      RECT 20.5000 1011.0850 119.5000 1012.3150 ;
      RECT 920.5700 1010.5150 999.5000 1011.0850 ;
      RECT 900.5000 1010.5150 920.0000 1011.0850 ;
      RECT 99.8350 1010.5150 119.5000 1011.0850 ;
      RECT 20.5000 1010.5150 99.2650 1011.0850 ;
      RECT 900.5000 1009.2850 999.5000 1010.5150 ;
      RECT 20.5000 1009.2850 119.5000 1010.5150 ;
      RECT 920.5700 1008.7150 999.5000 1009.2850 ;
      RECT 900.5000 1008.7150 920.0000 1009.2850 ;
      RECT 99.8350 1008.7150 119.5000 1009.2850 ;
      RECT 20.5000 1008.7150 99.2650 1009.2850 ;
      RECT 900.5000 1007.4850 999.5000 1008.7150 ;
      RECT 20.5000 1007.4850 119.5000 1008.7150 ;
      RECT 920.5700 1006.9150 999.5000 1007.4850 ;
      RECT 900.5000 1006.9150 920.0000 1007.4850 ;
      RECT 99.8350 1006.9150 119.5000 1007.4850 ;
      RECT 20.5000 1006.9150 99.2650 1007.4850 ;
      RECT 900.5000 1005.6850 999.5000 1006.9150 ;
      RECT 20.5000 1005.6850 119.5000 1006.9150 ;
      RECT 920.5700 1005.1150 999.5000 1005.6850 ;
      RECT 900.5000 1005.1150 920.0000 1005.6850 ;
      RECT 99.8350 1005.1150 119.5000 1005.6850 ;
      RECT 20.5000 1005.1150 99.2650 1005.6850 ;
      RECT 900.5000 1003.8850 999.5000 1005.1150 ;
      RECT 20.5000 1003.8850 119.5000 1005.1150 ;
      RECT 920.5700 1003.3150 999.5000 1003.8850 ;
      RECT 900.5000 1003.3150 920.0000 1003.8850 ;
      RECT 99.8350 1003.3150 119.5000 1003.8850 ;
      RECT 20.5000 1003.3150 99.2650 1003.8850 ;
      RECT 900.5000 1002.0850 999.5000 1003.3150 ;
      RECT 20.5000 1002.0850 119.5000 1003.3150 ;
      RECT 920.5700 1001.5150 999.5000 1002.0850 ;
      RECT 900.5000 1001.5150 920.0000 1002.0850 ;
      RECT 99.8350 1001.5150 119.5000 1002.0850 ;
      RECT 20.5000 1001.5150 99.2650 1002.0850 ;
      RECT 900.5000 1000.2850 999.5000 1001.5150 ;
      RECT 20.5000 1000.2850 119.5000 1001.5150 ;
      RECT 920.5700 999.7150 999.5000 1000.2850 ;
      RECT 900.5000 999.7150 920.0000 1000.2850 ;
      RECT 99.8350 999.7150 119.5000 1000.2850 ;
      RECT 20.5000 999.7150 99.2650 1000.2850 ;
      RECT 900.5000 998.4850 999.5000 999.7150 ;
      RECT 20.5000 998.4850 119.5000 999.7150 ;
      RECT 920.5700 997.9150 999.5000 998.4850 ;
      RECT 900.5000 997.9150 920.0000 998.4850 ;
      RECT 99.8350 997.9150 119.5000 998.4850 ;
      RECT 20.5000 997.9150 99.2650 998.4850 ;
      RECT 900.5000 996.6850 999.5000 997.9150 ;
      RECT 20.5000 996.6850 119.5000 997.9150 ;
      RECT 920.5700 996.1150 999.5000 996.6850 ;
      RECT 900.5000 996.1150 920.0000 996.6850 ;
      RECT 99.8350 996.1150 119.5000 996.6850 ;
      RECT 20.5000 996.1150 99.2650 996.6850 ;
      RECT 900.5000 994.8850 999.5000 996.1150 ;
      RECT 20.5000 994.8850 119.5000 996.1150 ;
      RECT 920.5700 994.3150 999.5000 994.8850 ;
      RECT 900.5000 994.3150 920.0000 994.8850 ;
      RECT 99.8350 994.3150 119.5000 994.8850 ;
      RECT 20.5000 994.3150 99.2650 994.8850 ;
      RECT 900.5000 993.0850 999.5000 994.3150 ;
      RECT 20.5000 993.0850 119.5000 994.3150 ;
      RECT 920.5700 992.5150 999.5000 993.0850 ;
      RECT 900.5000 992.5150 920.0000 993.0850 ;
      RECT 99.8350 992.5150 119.5000 993.0850 ;
      RECT 20.5000 992.5150 99.2650 993.0850 ;
      RECT 900.5000 991.2850 999.5000 992.5150 ;
      RECT 20.5000 991.2850 119.5000 992.5150 ;
      RECT 920.5700 990.7150 999.5000 991.2850 ;
      RECT 900.5000 990.7150 920.0000 991.2850 ;
      RECT 99.8350 990.7150 119.5000 991.2850 ;
      RECT 20.5000 990.7150 99.2650 991.2850 ;
      RECT 900.5000 989.4850 999.5000 990.7150 ;
      RECT 20.5000 989.4850 119.5000 990.7150 ;
      RECT 920.5700 988.9150 999.5000 989.4850 ;
      RECT 900.5000 988.9150 920.0000 989.4850 ;
      RECT 99.8350 988.9150 119.5000 989.4850 ;
      RECT 20.5000 988.9150 99.2650 989.4850 ;
      RECT 900.5000 987.6850 999.5000 988.9150 ;
      RECT 20.5000 987.6850 119.5000 988.9150 ;
      RECT 920.5700 987.1150 999.5000 987.6850 ;
      RECT 900.5000 987.1150 920.0000 987.6850 ;
      RECT 99.8350 987.1150 119.5000 987.6850 ;
      RECT 20.5000 987.1150 99.2650 987.6850 ;
      RECT 900.5000 985.8850 999.5000 987.1150 ;
      RECT 20.5000 985.8850 119.5000 987.1150 ;
      RECT 920.5700 985.3150 999.5000 985.8850 ;
      RECT 900.5000 985.3150 920.0000 985.8850 ;
      RECT 99.8350 985.3150 119.5000 985.8850 ;
      RECT 20.5000 985.3150 99.2650 985.8850 ;
      RECT 900.5000 984.0850 999.5000 985.3150 ;
      RECT 20.5000 984.0850 119.5000 985.3150 ;
      RECT 920.5700 983.5150 999.5000 984.0850 ;
      RECT 900.5000 983.5150 920.0000 984.0850 ;
      RECT 99.8350 983.5150 119.5000 984.0850 ;
      RECT 20.5000 983.5150 99.2650 984.0850 ;
      RECT 900.5000 982.2850 999.5000 983.5150 ;
      RECT 20.5000 982.2850 119.5000 983.5150 ;
      RECT 920.5700 981.7150 999.5000 982.2850 ;
      RECT 900.5000 981.7150 920.0000 982.2850 ;
      RECT 99.8350 981.7150 119.5000 982.2850 ;
      RECT 20.5000 981.7150 99.2650 982.2850 ;
      RECT 900.5000 980.4850 999.5000 981.7150 ;
      RECT 20.5000 980.4850 119.5000 981.7150 ;
      RECT 920.5700 979.9150 999.5000 980.4850 ;
      RECT 900.5000 979.9150 920.0000 980.4850 ;
      RECT 99.8350 979.9150 119.5000 980.4850 ;
      RECT 20.5000 979.9150 99.2650 980.4850 ;
      RECT 900.5000 978.6850 999.5000 979.9150 ;
      RECT 20.5000 978.6850 119.5000 979.9150 ;
      RECT 920.5700 978.1150 999.5000 978.6850 ;
      RECT 900.5000 978.1150 920.0000 978.6850 ;
      RECT 99.8350 978.1150 119.5000 978.6850 ;
      RECT 20.5000 978.1150 99.2650 978.6850 ;
      RECT 900.5000 976.8850 999.5000 978.1150 ;
      RECT 20.5000 976.8850 119.5000 978.1150 ;
      RECT 920.5700 976.3150 999.5000 976.8850 ;
      RECT 900.5000 976.3150 920.0000 976.8850 ;
      RECT 99.8350 976.3150 119.5000 976.8850 ;
      RECT 20.5000 976.3150 99.2650 976.8850 ;
      RECT 900.5000 975.0850 999.5000 976.3150 ;
      RECT 20.5000 975.0850 119.5000 976.3150 ;
      RECT 920.5700 974.5150 999.5000 975.0850 ;
      RECT 900.5000 974.5150 920.0000 975.0850 ;
      RECT 99.8350 974.5150 119.5000 975.0850 ;
      RECT 20.5000 974.5150 99.2650 975.0850 ;
      RECT 900.5000 973.2850 999.5000 974.5150 ;
      RECT 20.5000 973.2850 119.5000 974.5150 ;
      RECT 920.5700 972.7150 999.5000 973.2850 ;
      RECT 900.5000 972.7150 920.0000 973.2850 ;
      RECT 99.8350 972.7150 119.5000 973.2850 ;
      RECT 20.5000 972.7150 99.2650 973.2850 ;
      RECT 900.5000 971.4850 999.5000 972.7150 ;
      RECT 20.5000 971.4850 119.5000 972.7150 ;
      RECT 920.5700 970.9150 999.5000 971.4850 ;
      RECT 900.5000 970.9150 920.0000 971.4850 ;
      RECT 99.8350 970.9150 119.5000 971.4850 ;
      RECT 20.5000 970.9150 99.2650 971.4850 ;
      RECT 900.5000 969.6850 999.5000 970.9150 ;
      RECT 20.5000 969.6850 119.5000 970.9150 ;
      RECT 920.5700 969.1150 999.5000 969.6850 ;
      RECT 900.5000 969.1150 920.0000 969.6850 ;
      RECT 99.8350 969.1150 119.5000 969.6850 ;
      RECT 20.5000 969.1150 99.2650 969.6850 ;
      RECT 900.5000 967.8850 999.5000 969.1150 ;
      RECT 20.5000 967.8850 119.5000 969.1150 ;
      RECT 920.5700 967.3150 999.5000 967.8850 ;
      RECT 900.5000 967.3150 920.0000 967.8850 ;
      RECT 99.8350 967.3150 119.5000 967.8850 ;
      RECT 20.5000 967.3150 99.2650 967.8850 ;
      RECT 900.5000 966.0850 999.5000 967.3150 ;
      RECT 20.5000 966.0850 119.5000 967.3150 ;
      RECT 920.5700 965.5150 999.5000 966.0850 ;
      RECT 900.5000 965.5150 920.0000 966.0850 ;
      RECT 99.8350 965.5150 119.5000 966.0850 ;
      RECT 20.5000 965.5150 99.2650 966.0850 ;
      RECT 900.5000 964.2850 999.5000 965.5150 ;
      RECT 20.5000 964.2850 119.5000 965.5150 ;
      RECT 920.5700 963.7150 999.5000 964.2850 ;
      RECT 900.5000 963.7150 920.0000 964.2850 ;
      RECT 99.8350 963.7150 119.5000 964.2850 ;
      RECT 20.5000 963.7150 99.2650 964.2850 ;
      RECT 900.5000 962.4850 999.5000 963.7150 ;
      RECT 20.5000 962.4850 119.5000 963.7150 ;
      RECT 920.5700 961.9150 999.5000 962.4850 ;
      RECT 900.5000 961.9150 920.0000 962.4850 ;
      RECT 99.8350 961.9150 119.5000 962.4850 ;
      RECT 20.5000 961.9150 99.2650 962.4850 ;
      RECT 900.5000 960.6850 999.5000 961.9150 ;
      RECT 20.5000 960.6850 119.5000 961.9150 ;
      RECT 920.5700 960.1150 999.5000 960.6850 ;
      RECT 900.5000 960.1150 920.0000 960.6850 ;
      RECT 99.8350 960.1150 119.5000 960.6850 ;
      RECT 20.5000 960.1150 99.2650 960.6850 ;
      RECT 900.5000 958.8850 999.5000 960.1150 ;
      RECT 20.5000 958.8850 119.5000 960.1150 ;
      RECT 920.5700 958.3150 999.5000 958.8850 ;
      RECT 900.5000 958.3150 920.0000 958.8850 ;
      RECT 99.8350 958.3150 119.5000 958.8850 ;
      RECT 20.5000 958.3150 99.2650 958.8850 ;
      RECT 900.5000 957.0850 999.5000 958.3150 ;
      RECT 20.5000 957.0850 119.5000 958.3150 ;
      RECT 920.5700 956.5150 999.5000 957.0850 ;
      RECT 900.5000 956.5150 920.0000 957.0850 ;
      RECT 99.8350 956.5150 119.5000 957.0850 ;
      RECT 20.5000 956.5150 99.2650 957.0850 ;
      RECT 900.5000 955.2850 999.5000 956.5150 ;
      RECT 20.5000 955.2850 119.5000 956.5150 ;
      RECT 920.5700 954.7150 999.5000 955.2850 ;
      RECT 900.5000 954.7150 920.0000 955.2850 ;
      RECT 99.8350 954.7150 119.5000 955.2850 ;
      RECT 20.5000 954.7150 99.2650 955.2850 ;
      RECT 900.5000 953.4850 999.5000 954.7150 ;
      RECT 20.5000 953.4850 119.5000 954.7150 ;
      RECT 920.5700 952.9150 999.5000 953.4850 ;
      RECT 900.5000 952.9150 920.0000 953.4850 ;
      RECT 99.8350 952.9150 119.5000 953.4850 ;
      RECT 20.5000 952.9150 99.2650 953.4850 ;
      RECT 900.5000 951.6850 999.5000 952.9150 ;
      RECT 20.5000 951.6850 119.5000 952.9150 ;
      RECT 920.5700 951.1150 999.5000 951.6850 ;
      RECT 900.5000 951.1150 920.0000 951.6850 ;
      RECT 99.8350 951.1150 119.5000 951.6850 ;
      RECT 20.5000 951.1150 99.2650 951.6850 ;
      RECT 900.5000 949.8850 999.5000 951.1150 ;
      RECT 20.5000 949.8850 119.5000 951.1150 ;
      RECT 920.5700 949.3150 999.5000 949.8850 ;
      RECT 900.5000 949.3150 920.0000 949.8850 ;
      RECT 99.8350 949.3150 119.5000 949.8850 ;
      RECT 20.5000 949.3150 99.2650 949.8850 ;
      RECT 900.5000 948.0850 999.5000 949.3150 ;
      RECT 20.5000 948.0850 119.5000 949.3150 ;
      RECT 920.5700 947.5150 999.5000 948.0850 ;
      RECT 900.5000 947.5150 920.0000 948.0850 ;
      RECT 99.8350 947.5150 119.5000 948.0850 ;
      RECT 20.5000 947.5150 99.2650 948.0850 ;
      RECT 900.5000 946.2850 999.5000 947.5150 ;
      RECT 20.5000 946.2850 119.5000 947.5150 ;
      RECT 920.5700 945.7150 999.5000 946.2850 ;
      RECT 900.5000 945.7150 920.0000 946.2850 ;
      RECT 99.8350 945.7150 119.5000 946.2850 ;
      RECT 20.5000 945.7150 99.2650 946.2850 ;
      RECT 900.5000 944.4850 999.5000 945.7150 ;
      RECT 20.5000 944.4850 119.5000 945.7150 ;
      RECT 920.5700 943.9150 999.5000 944.4850 ;
      RECT 900.5000 943.9150 920.0000 944.4850 ;
      RECT 99.8350 943.9150 119.5000 944.4850 ;
      RECT 20.5000 943.9150 99.2650 944.4850 ;
      RECT 900.5000 942.6850 999.5000 943.9150 ;
      RECT 20.5000 942.6850 119.5000 943.9150 ;
      RECT 920.5700 942.1150 999.5000 942.6850 ;
      RECT 900.5000 942.1150 920.0000 942.6850 ;
      RECT 99.8350 942.1150 119.5000 942.6850 ;
      RECT 20.5000 942.1150 99.2650 942.6850 ;
      RECT 900.5000 940.8850 999.5000 942.1150 ;
      RECT 20.5000 940.8850 119.5000 942.1150 ;
      RECT 920.5700 940.3150 999.5000 940.8850 ;
      RECT 900.5000 940.3150 920.0000 940.8850 ;
      RECT 99.8350 940.3150 119.5000 940.8850 ;
      RECT 20.5000 940.3150 99.2650 940.8850 ;
      RECT 900.5000 939.0850 999.5000 940.3150 ;
      RECT 20.5000 939.0850 119.5000 940.3150 ;
      RECT 920.5700 938.5150 999.5000 939.0850 ;
      RECT 900.5000 938.5150 920.0000 939.0850 ;
      RECT 99.8350 938.5150 119.5000 939.0850 ;
      RECT 20.5000 938.5150 99.2650 939.0850 ;
      RECT 900.5000 937.2850 999.5000 938.5150 ;
      RECT 20.5000 937.2850 119.5000 938.5150 ;
      RECT 920.5700 936.7150 999.5000 937.2850 ;
      RECT 900.5000 936.7150 920.0000 937.2850 ;
      RECT 99.8350 936.7150 119.5000 937.2850 ;
      RECT 20.5000 936.7150 99.2650 937.2850 ;
      RECT 900.5000 935.4850 999.5000 936.7150 ;
      RECT 20.5000 935.4850 119.5000 936.7150 ;
      RECT 920.5700 934.9150 999.5000 935.4850 ;
      RECT 900.5000 934.9150 920.0000 935.4850 ;
      RECT 99.8350 934.9150 119.5000 935.4850 ;
      RECT 20.5000 934.9150 99.2650 935.4850 ;
      RECT 900.5000 933.6850 999.5000 934.9150 ;
      RECT 20.5000 933.6850 119.5000 934.9150 ;
      RECT 920.5700 933.1150 999.5000 933.6850 ;
      RECT 900.5000 933.1150 920.0000 933.6850 ;
      RECT 99.8350 933.1150 119.5000 933.6850 ;
      RECT 20.5000 933.1150 99.2650 933.6850 ;
      RECT 900.5000 931.8850 999.5000 933.1150 ;
      RECT 20.5000 931.8850 119.5000 933.1150 ;
      RECT 920.5700 931.3150 999.5000 931.8850 ;
      RECT 900.5000 931.3150 920.0000 931.8850 ;
      RECT 99.8350 931.3150 119.5000 931.8850 ;
      RECT 20.5000 931.3150 99.2650 931.8850 ;
      RECT 900.5000 930.0850 999.5000 931.3150 ;
      RECT 20.5000 930.0850 119.5000 931.3150 ;
      RECT 920.5700 929.5150 999.5000 930.0850 ;
      RECT 900.5000 929.5150 920.0000 930.0850 ;
      RECT 99.8350 929.5150 119.5000 930.0850 ;
      RECT 20.5000 929.5150 99.2650 930.0850 ;
      RECT 900.5000 928.2850 999.5000 929.5150 ;
      RECT 20.5000 928.2850 119.5000 929.5150 ;
      RECT 920.5700 927.7150 999.5000 928.2850 ;
      RECT 900.5000 927.7150 920.0000 928.2850 ;
      RECT 99.8350 927.7150 119.5000 928.2850 ;
      RECT 20.5000 927.7150 99.2650 928.2850 ;
      RECT 900.5000 926.4850 999.5000 927.7150 ;
      RECT 20.5000 926.4850 119.5000 927.7150 ;
      RECT 920.5700 925.9150 999.5000 926.4850 ;
      RECT 900.5000 925.9150 920.0000 926.4850 ;
      RECT 99.8350 925.9150 119.5000 926.4850 ;
      RECT 20.5000 925.9150 99.2650 926.4850 ;
      RECT 900.5000 924.6850 999.5000 925.9150 ;
      RECT 20.5000 924.6850 119.5000 925.9150 ;
      RECT 920.5700 924.1150 999.5000 924.6850 ;
      RECT 900.5000 924.1150 920.0000 924.6850 ;
      RECT 99.8350 924.1150 119.5000 924.6850 ;
      RECT 20.5000 924.1150 99.2650 924.6850 ;
      RECT 900.5000 922.8850 999.5000 924.1150 ;
      RECT 20.5000 922.8850 119.5000 924.1150 ;
      RECT 920.5700 922.3150 999.5000 922.8850 ;
      RECT 900.5000 922.3150 920.0000 922.8850 ;
      RECT 99.8350 922.3150 119.5000 922.8850 ;
      RECT 20.5000 922.3150 99.2650 922.8850 ;
      RECT 900.5000 921.0850 999.5000 922.3150 ;
      RECT 20.5000 921.0850 119.5000 922.3150 ;
      RECT 920.5700 920.5150 999.5000 921.0850 ;
      RECT 900.5000 920.5150 920.0000 921.0850 ;
      RECT 99.8350 920.5150 119.5000 921.0850 ;
      RECT 20.5000 920.5150 99.2650 921.0850 ;
      RECT 900.5000 919.2850 999.5000 920.5150 ;
      RECT 20.5000 919.2850 119.5000 920.5150 ;
      RECT 920.5700 918.7150 999.5000 919.2850 ;
      RECT 900.5000 918.7150 920.0000 919.2850 ;
      RECT 99.8350 918.7150 119.5000 919.2850 ;
      RECT 20.5000 918.7150 99.2650 919.2850 ;
      RECT 900.5000 917.4850 999.5000 918.7150 ;
      RECT 20.5000 917.4850 119.5000 918.7150 ;
      RECT 920.5700 916.9150 999.5000 917.4850 ;
      RECT 900.5000 916.9150 920.0000 917.4850 ;
      RECT 99.8350 916.9150 119.5000 917.4850 ;
      RECT 20.5000 916.9150 99.2650 917.4850 ;
      RECT 900.5000 915.6850 999.5000 916.9150 ;
      RECT 20.5000 915.6850 119.5000 916.9150 ;
      RECT 920.5700 915.1150 999.5000 915.6850 ;
      RECT 900.5000 915.1150 920.0000 915.6850 ;
      RECT 99.8350 915.1150 119.5000 915.6850 ;
      RECT 20.5000 915.1150 99.2650 915.6850 ;
      RECT 900.5000 913.8850 999.5000 915.1150 ;
      RECT 20.5000 913.8850 119.5000 915.1150 ;
      RECT 920.5700 913.3150 999.5000 913.8850 ;
      RECT 900.5000 913.3150 920.0000 913.8850 ;
      RECT 99.8350 913.3150 119.5000 913.8850 ;
      RECT 20.5000 913.3150 99.2650 913.8850 ;
      RECT 900.5000 912.0850 999.5000 913.3150 ;
      RECT 20.5000 912.0850 119.5000 913.3150 ;
      RECT 920.5700 911.5150 999.5000 912.0850 ;
      RECT 900.5000 911.5150 920.0000 912.0850 ;
      RECT 99.8350 911.5150 119.5000 912.0850 ;
      RECT 20.5000 911.5150 99.2650 912.0850 ;
      RECT 900.5000 910.2850 999.5000 911.5150 ;
      RECT 20.5000 910.2850 119.5000 911.5150 ;
      RECT 920.5700 909.7150 999.5000 910.2850 ;
      RECT 900.5000 909.7150 920.0000 910.2850 ;
      RECT 99.8350 909.7150 119.5000 910.2850 ;
      RECT 20.5000 909.7150 99.2650 910.2850 ;
      RECT 900.5000 908.4850 999.5000 909.7150 ;
      RECT 20.5000 908.4850 119.5000 909.7150 ;
      RECT 920.5700 907.9150 999.5000 908.4850 ;
      RECT 900.5000 907.9150 920.0000 908.4850 ;
      RECT 99.8350 907.9150 119.5000 908.4850 ;
      RECT 20.5000 907.9150 99.2650 908.4850 ;
      RECT 900.5000 906.6850 999.5000 907.9150 ;
      RECT 20.5000 906.6850 119.5000 907.9150 ;
      RECT 920.5700 906.1150 999.5000 906.6850 ;
      RECT 900.5000 906.1150 920.0000 906.6850 ;
      RECT 99.8350 906.1150 119.5000 906.6850 ;
      RECT 20.5000 906.1150 99.2650 906.6850 ;
      RECT 900.5000 904.8850 999.5000 906.1150 ;
      RECT 20.5000 904.8850 119.5000 906.1150 ;
      RECT 920.5700 904.3150 999.5000 904.8850 ;
      RECT 900.5000 904.3150 920.0000 904.8850 ;
      RECT 99.8350 904.3150 119.5000 904.8850 ;
      RECT 20.5000 904.3150 99.2650 904.8850 ;
      RECT 900.5000 903.0850 999.5000 904.3150 ;
      RECT 20.5000 903.0850 119.5000 904.3150 ;
      RECT 920.5700 902.5150 999.5000 903.0850 ;
      RECT 900.5000 902.5150 920.0000 903.0850 ;
      RECT 99.8350 902.5150 119.5000 903.0850 ;
      RECT 20.5000 902.5150 99.2650 903.0850 ;
      RECT 900.5000 901.2850 999.5000 902.5150 ;
      RECT 20.5000 901.2850 119.5000 902.5150 ;
      RECT 920.5700 900.7150 999.5000 901.2850 ;
      RECT 900.5000 900.7150 920.0000 901.2850 ;
      RECT 99.8350 900.7150 119.5000 901.2850 ;
      RECT 20.5000 900.7150 99.2650 901.2850 ;
      RECT 900.5000 899.4850 999.5000 900.7150 ;
      RECT 20.5000 899.4850 119.5000 900.7150 ;
      RECT 920.5700 898.9150 999.5000 899.4850 ;
      RECT 900.5000 898.9150 920.0000 899.4850 ;
      RECT 99.8350 898.9150 119.5000 899.4850 ;
      RECT 20.5000 898.9150 99.2650 899.4850 ;
      RECT 900.5000 897.6850 999.5000 898.9150 ;
      RECT 20.5000 897.6850 119.5000 898.9150 ;
      RECT 920.5700 897.1150 999.5000 897.6850 ;
      RECT 900.5000 897.1150 920.0000 897.6850 ;
      RECT 99.8350 897.1150 119.5000 897.6850 ;
      RECT 20.5000 897.1150 99.2650 897.6850 ;
      RECT 900.5000 895.8850 999.5000 897.1150 ;
      RECT 20.5000 895.8850 119.5000 897.1150 ;
      RECT 920.5700 895.3150 999.5000 895.8850 ;
      RECT 900.5000 895.3150 920.0000 895.8850 ;
      RECT 99.8350 895.3150 119.5000 895.8850 ;
      RECT 20.5000 895.3150 99.2650 895.8850 ;
      RECT 900.5000 894.0850 999.5000 895.3150 ;
      RECT 20.5000 894.0850 119.5000 895.3150 ;
      RECT 920.5700 893.5150 999.5000 894.0850 ;
      RECT 900.5000 893.5150 920.0000 894.0850 ;
      RECT 99.8350 893.5150 119.5000 894.0850 ;
      RECT 20.5000 893.5150 99.2650 894.0850 ;
      RECT 900.5000 892.2850 999.5000 893.5150 ;
      RECT 20.5000 892.2850 119.5000 893.5150 ;
      RECT 920.5700 891.7150 999.5000 892.2850 ;
      RECT 900.5000 891.7150 920.0000 892.2850 ;
      RECT 99.8350 891.7150 119.5000 892.2850 ;
      RECT 20.5000 891.7150 99.2650 892.2850 ;
      RECT 900.5000 890.4850 999.5000 891.7150 ;
      RECT 20.5000 890.4850 119.5000 891.7150 ;
      RECT 920.5700 889.9150 999.5000 890.4850 ;
      RECT 900.5000 889.9150 920.0000 890.4850 ;
      RECT 99.8350 889.9150 119.5000 890.4850 ;
      RECT 20.5000 889.9150 99.2650 890.4850 ;
      RECT 900.5000 888.6850 999.5000 889.9150 ;
      RECT 20.5000 888.6850 119.5000 889.9150 ;
      RECT 920.5700 888.1150 999.5000 888.6850 ;
      RECT 900.5000 888.1150 920.0000 888.6850 ;
      RECT 99.8350 888.1150 119.5000 888.6850 ;
      RECT 20.5000 888.1150 99.2650 888.6850 ;
      RECT 900.5000 886.8850 999.5000 888.1150 ;
      RECT 20.5000 886.8850 119.5000 888.1150 ;
      RECT 920.5700 886.3150 999.5000 886.8850 ;
      RECT 900.5000 886.3150 920.0000 886.8850 ;
      RECT 99.8350 886.3150 119.5000 886.8850 ;
      RECT 20.5000 886.3150 99.2650 886.8850 ;
      RECT 900.5000 885.0850 999.5000 886.3150 ;
      RECT 20.5000 885.0850 119.5000 886.3150 ;
      RECT 920.5700 884.5150 999.5000 885.0850 ;
      RECT 900.5000 884.5150 920.0000 885.0850 ;
      RECT 99.8350 884.5150 119.5000 885.0850 ;
      RECT 20.5000 884.5150 99.2650 885.0850 ;
      RECT 900.5000 883.2850 999.5000 884.5150 ;
      RECT 20.5000 883.2850 119.5000 884.5150 ;
      RECT 920.5700 882.7150 999.5000 883.2850 ;
      RECT 900.5000 882.7150 920.0000 883.2850 ;
      RECT 99.8350 882.7150 119.5000 883.2850 ;
      RECT 20.5000 882.7150 99.2650 883.2850 ;
      RECT 900.5000 881.4850 999.5000 882.7150 ;
      RECT 20.5000 881.4850 119.5000 882.7150 ;
      RECT 920.5700 880.9150 999.5000 881.4850 ;
      RECT 900.5000 880.9150 920.0000 881.4850 ;
      RECT 99.8350 880.9150 119.5000 881.4850 ;
      RECT 20.5000 880.9150 99.2650 881.4850 ;
      RECT 900.5000 879.6850 999.5000 880.9150 ;
      RECT 20.5000 879.6850 119.5000 880.9150 ;
      RECT 920.5700 879.1150 999.5000 879.6850 ;
      RECT 900.5000 879.1150 920.0000 879.6850 ;
      RECT 99.8350 879.1150 119.5000 879.6850 ;
      RECT 20.5000 879.1150 99.2650 879.6850 ;
      RECT 900.5000 877.8850 999.5000 879.1150 ;
      RECT 20.5000 877.8850 119.5000 879.1150 ;
      RECT 920.5700 877.3150 999.5000 877.8850 ;
      RECT 900.5000 877.3150 920.0000 877.8850 ;
      RECT 99.8350 877.3150 119.5000 877.8850 ;
      RECT 20.5000 877.3150 99.2650 877.8850 ;
      RECT 900.5000 876.0850 999.5000 877.3150 ;
      RECT 20.5000 876.0850 119.5000 877.3150 ;
      RECT 920.5700 875.5150 999.5000 876.0850 ;
      RECT 900.5000 875.5150 920.0000 876.0850 ;
      RECT 99.8350 875.5150 119.5000 876.0850 ;
      RECT 20.5000 875.5150 99.2650 876.0850 ;
      RECT 900.5000 874.2850 999.5000 875.5150 ;
      RECT 20.5000 874.2850 119.5000 875.5150 ;
      RECT 920.5700 873.7150 999.5000 874.2850 ;
      RECT 900.5000 873.7150 920.0000 874.2850 ;
      RECT 99.8350 873.7150 119.5000 874.2850 ;
      RECT 20.5000 873.7150 99.2650 874.2850 ;
      RECT 900.5000 872.4850 999.5000 873.7150 ;
      RECT 20.5000 872.4850 119.5000 873.7150 ;
      RECT 920.5700 871.9150 999.5000 872.4850 ;
      RECT 900.5000 871.9150 920.0000 872.4850 ;
      RECT 99.8350 871.9150 119.5000 872.4850 ;
      RECT 20.5000 871.9150 99.2650 872.4850 ;
      RECT 900.5000 870.6850 999.5000 871.9150 ;
      RECT 20.5000 870.6850 119.5000 871.9150 ;
      RECT 920.5700 870.1150 999.5000 870.6850 ;
      RECT 900.5000 870.1150 920.0000 870.6850 ;
      RECT 99.8350 870.1150 119.5000 870.6850 ;
      RECT 20.5000 870.1150 99.2650 870.6850 ;
      RECT 900.5000 868.8850 999.5000 870.1150 ;
      RECT 20.5000 868.8850 119.5000 870.1150 ;
      RECT 920.5700 868.3150 999.5000 868.8850 ;
      RECT 900.5000 868.3150 920.0000 868.8850 ;
      RECT 99.8350 868.3150 119.5000 868.8850 ;
      RECT 20.5000 868.3150 99.2650 868.8850 ;
      RECT 900.5000 867.0850 999.5000 868.3150 ;
      RECT 20.5000 867.0850 119.5000 868.3150 ;
      RECT 920.5700 866.5150 999.5000 867.0850 ;
      RECT 900.5000 866.5150 920.0000 867.0850 ;
      RECT 99.8350 866.5150 119.5000 867.0850 ;
      RECT 20.5000 866.5150 99.2650 867.0850 ;
      RECT 900.5000 865.2850 999.5000 866.5150 ;
      RECT 20.5000 865.2850 119.5000 866.5150 ;
      RECT 920.5700 864.7150 999.5000 865.2850 ;
      RECT 900.5000 864.7150 920.0000 865.2850 ;
      RECT 99.8350 864.7150 119.5000 865.2850 ;
      RECT 20.5000 864.7150 99.2650 865.2850 ;
      RECT 900.5000 863.4850 999.5000 864.7150 ;
      RECT 20.5000 863.4850 119.5000 864.7150 ;
      RECT 920.5700 862.9150 999.5000 863.4850 ;
      RECT 900.5000 862.9150 920.0000 863.4850 ;
      RECT 99.8350 862.9150 119.5000 863.4850 ;
      RECT 20.5000 862.9150 99.2650 863.4850 ;
      RECT 900.5000 861.6850 999.5000 862.9150 ;
      RECT 20.5000 861.6850 119.5000 862.9150 ;
      RECT 920.5700 861.1150 999.5000 861.6850 ;
      RECT 900.5000 861.1150 920.0000 861.6850 ;
      RECT 99.8350 861.1150 119.5000 861.6850 ;
      RECT 20.5000 861.1150 99.2650 861.6850 ;
      RECT 900.5000 859.8850 999.5000 861.1150 ;
      RECT 20.5000 859.8850 119.5000 861.1150 ;
      RECT 920.5700 859.3150 999.5000 859.8850 ;
      RECT 900.5000 859.3150 920.0000 859.8850 ;
      RECT 99.8350 859.3150 119.5000 859.8850 ;
      RECT 20.5000 859.3150 99.2650 859.8850 ;
      RECT 900.5000 858.0850 999.5000 859.3150 ;
      RECT 20.5000 858.0850 119.5000 859.3150 ;
      RECT 920.5700 857.5150 999.5000 858.0850 ;
      RECT 900.5000 857.5150 920.0000 858.0850 ;
      RECT 99.8350 857.5150 119.5000 858.0850 ;
      RECT 20.5000 857.5150 99.2650 858.0850 ;
      RECT 900.5000 856.2850 999.5000 857.5150 ;
      RECT 20.5000 856.2850 119.5000 857.5150 ;
      RECT 920.5700 855.7150 999.5000 856.2850 ;
      RECT 900.5000 855.7150 920.0000 856.2850 ;
      RECT 99.8350 855.7150 119.5000 856.2850 ;
      RECT 20.5000 855.7150 99.2650 856.2850 ;
      RECT 900.5000 854.4850 999.5000 855.7150 ;
      RECT 20.5000 854.4850 119.5000 855.7150 ;
      RECT 920.5700 853.9150 999.5000 854.4850 ;
      RECT 900.5000 853.9150 920.0000 854.4850 ;
      RECT 99.8350 853.9150 119.5000 854.4850 ;
      RECT 20.5000 853.9150 99.2650 854.4850 ;
      RECT 900.5000 852.6850 999.5000 853.9150 ;
      RECT 20.5000 852.6850 119.5000 853.9150 ;
      RECT 920.5700 852.1150 999.5000 852.6850 ;
      RECT 900.5000 852.1150 920.0000 852.6850 ;
      RECT 99.8350 852.1150 119.5000 852.6850 ;
      RECT 20.5000 852.1150 99.2650 852.6850 ;
      RECT 900.5000 850.8850 999.5000 852.1150 ;
      RECT 20.5000 850.8850 119.5000 852.1150 ;
      RECT 920.5700 850.3150 999.5000 850.8850 ;
      RECT 900.5000 850.3150 920.0000 850.8850 ;
      RECT 99.8350 850.3150 119.5000 850.8850 ;
      RECT 20.5000 850.3150 99.2650 850.8850 ;
      RECT 900.5000 849.0850 999.5000 850.3150 ;
      RECT 20.5000 849.0850 119.5000 850.3150 ;
      RECT 920.5700 848.5150 999.5000 849.0850 ;
      RECT 900.5000 848.5150 920.0000 849.0850 ;
      RECT 99.8350 848.5150 119.5000 849.0850 ;
      RECT 20.5000 848.5150 99.2650 849.0850 ;
      RECT 900.5000 847.2850 999.5000 848.5150 ;
      RECT 20.5000 847.2850 119.5000 848.5150 ;
      RECT 920.5700 846.7150 999.5000 847.2850 ;
      RECT 900.5000 846.7150 920.0000 847.2850 ;
      RECT 99.8350 846.7150 119.5000 847.2850 ;
      RECT 20.5000 846.7150 99.2650 847.2850 ;
      RECT 900.5000 845.4850 999.5000 846.7150 ;
      RECT 20.5000 845.4850 119.5000 846.7150 ;
      RECT 920.5700 844.9150 999.5000 845.4850 ;
      RECT 900.5000 844.9150 920.0000 845.4850 ;
      RECT 99.8350 844.9150 119.5000 845.4850 ;
      RECT 20.5000 844.9150 99.2650 845.4850 ;
      RECT 900.5000 843.6850 999.5000 844.9150 ;
      RECT 20.5000 843.6850 119.5000 844.9150 ;
      RECT 920.5700 843.1150 999.5000 843.6850 ;
      RECT 900.5000 843.1150 920.0000 843.6850 ;
      RECT 99.8350 843.1150 119.5000 843.6850 ;
      RECT 20.5000 843.1150 99.2650 843.6850 ;
      RECT 900.5000 841.8850 999.5000 843.1150 ;
      RECT 20.5000 841.8850 119.5000 843.1150 ;
      RECT 920.5700 841.3150 999.5000 841.8850 ;
      RECT 900.5000 841.3150 920.0000 841.8850 ;
      RECT 99.8350 841.3150 119.5000 841.8850 ;
      RECT 20.5000 841.3150 99.2650 841.8850 ;
      RECT 900.5000 840.0850 999.5000 841.3150 ;
      RECT 20.5000 840.0850 119.5000 841.3150 ;
      RECT 920.5700 839.5150 999.5000 840.0850 ;
      RECT 900.5000 839.5150 920.0000 840.0850 ;
      RECT 99.8350 839.5150 119.5000 840.0850 ;
      RECT 20.5000 839.5150 99.2650 840.0850 ;
      RECT 900.5000 838.2850 999.5000 839.5150 ;
      RECT 20.5000 838.2850 119.5000 839.5150 ;
      RECT 920.5700 837.7150 999.5000 838.2850 ;
      RECT 900.5000 837.7150 920.0000 838.2850 ;
      RECT 99.8350 837.7150 119.5000 838.2850 ;
      RECT 20.5000 837.7150 99.2650 838.2850 ;
      RECT 900.5000 836.4850 999.5000 837.7150 ;
      RECT 20.5000 836.4850 119.5000 837.7150 ;
      RECT 920.5700 835.9150 999.5000 836.4850 ;
      RECT 900.5000 835.9150 920.0000 836.4850 ;
      RECT 99.8350 835.9150 119.5000 836.4850 ;
      RECT 20.5000 835.9150 99.2650 836.4850 ;
      RECT 900.5000 834.6850 999.5000 835.9150 ;
      RECT 20.5000 834.6850 119.5000 835.9150 ;
      RECT 920.5700 834.1150 999.5000 834.6850 ;
      RECT 900.5000 834.1150 920.0000 834.6850 ;
      RECT 99.8350 834.1150 119.5000 834.6850 ;
      RECT 20.5000 834.1150 99.2650 834.6850 ;
      RECT 900.5000 832.8850 999.5000 834.1150 ;
      RECT 20.5000 832.8850 119.5000 834.1150 ;
      RECT 920.5700 832.3150 999.5000 832.8850 ;
      RECT 900.5000 832.3150 920.0000 832.8850 ;
      RECT 99.8350 832.3150 119.5000 832.8850 ;
      RECT 20.5000 832.3150 99.2650 832.8850 ;
      RECT 900.5000 831.0850 999.5000 832.3150 ;
      RECT 20.5000 831.0850 119.5000 832.3150 ;
      RECT 920.5700 830.5150 999.5000 831.0850 ;
      RECT 900.5000 830.5150 920.0000 831.0850 ;
      RECT 99.8350 830.5150 119.5000 831.0850 ;
      RECT 20.5000 830.5150 99.2650 831.0850 ;
      RECT 900.5000 829.2850 999.5000 830.5150 ;
      RECT 20.5000 829.2850 119.5000 830.5150 ;
      RECT 920.5700 828.7150 999.5000 829.2850 ;
      RECT 900.5000 828.7150 920.0000 829.2850 ;
      RECT 99.8350 828.7150 119.5000 829.2850 ;
      RECT 20.5000 828.7150 99.2650 829.2850 ;
      RECT 900.5000 827.4850 999.5000 828.7150 ;
      RECT 20.5000 827.4850 119.5000 828.7150 ;
      RECT 920.5700 826.9150 999.5000 827.4850 ;
      RECT 900.5000 826.9150 920.0000 827.4850 ;
      RECT 99.8350 826.9150 119.5000 827.4850 ;
      RECT 20.5000 826.9150 99.2650 827.4850 ;
      RECT 900.5000 825.6850 999.5000 826.9150 ;
      RECT 20.5000 825.6850 119.5000 826.9150 ;
      RECT 920.5700 825.1150 999.5000 825.6850 ;
      RECT 900.5000 825.1150 920.0000 825.6850 ;
      RECT 99.8350 825.1150 119.5000 825.6850 ;
      RECT 20.5000 825.1150 99.2650 825.6850 ;
      RECT 900.5000 823.8850 999.5000 825.1150 ;
      RECT 20.5000 823.8850 119.5000 825.1150 ;
      RECT 920.5700 823.3150 999.5000 823.8850 ;
      RECT 900.5000 823.3150 920.0000 823.8850 ;
      RECT 99.8350 823.3150 119.5000 823.8850 ;
      RECT 20.5000 823.3150 99.2650 823.8850 ;
      RECT 900.5000 822.0850 999.5000 823.3150 ;
      RECT 20.5000 822.0850 119.5000 823.3150 ;
      RECT 920.5700 821.5150 999.5000 822.0850 ;
      RECT 900.5000 821.5150 920.0000 822.0850 ;
      RECT 99.8350 821.5150 119.5000 822.0850 ;
      RECT 20.5000 821.5150 99.2650 822.0850 ;
      RECT 900.5000 820.2850 999.5000 821.5150 ;
      RECT 20.5000 820.2850 119.5000 821.5150 ;
      RECT 920.5700 819.7150 999.5000 820.2850 ;
      RECT 900.5000 819.7150 920.0000 820.2850 ;
      RECT 99.8350 819.7150 119.5000 820.2850 ;
      RECT 20.5000 819.7150 99.2650 820.2850 ;
      RECT 900.5000 818.4850 999.5000 819.7150 ;
      RECT 20.5000 818.4850 119.5000 819.7150 ;
      RECT 920.5700 817.9150 999.5000 818.4850 ;
      RECT 900.5000 817.9150 920.0000 818.4850 ;
      RECT 99.8350 817.9150 119.5000 818.4850 ;
      RECT 20.5000 817.9150 99.2650 818.4850 ;
      RECT 900.5000 816.6850 999.5000 817.9150 ;
      RECT 20.5000 816.6850 119.5000 817.9150 ;
      RECT 920.5700 816.1150 999.5000 816.6850 ;
      RECT 900.5000 816.1150 920.0000 816.6850 ;
      RECT 99.8350 816.1150 119.5000 816.6850 ;
      RECT 20.5000 816.1150 99.2650 816.6850 ;
      RECT 900.5000 814.8850 999.5000 816.1150 ;
      RECT 20.5000 814.8850 119.5000 816.1150 ;
      RECT 920.5700 814.3150 999.5000 814.8850 ;
      RECT 900.5000 814.3150 920.0000 814.8850 ;
      RECT 99.8350 814.3150 119.5000 814.8850 ;
      RECT 20.5000 814.3150 99.2650 814.8850 ;
      RECT 900.5000 813.0850 999.5000 814.3150 ;
      RECT 20.5000 813.0850 119.5000 814.3150 ;
      RECT 920.5700 812.5150 999.5000 813.0850 ;
      RECT 900.5000 812.5150 920.0000 813.0850 ;
      RECT 99.8350 812.5150 119.5000 813.0850 ;
      RECT 20.5000 812.5150 99.2650 813.0850 ;
      RECT 900.5000 811.2850 999.5000 812.5150 ;
      RECT 20.5000 811.2850 119.5000 812.5150 ;
      RECT 920.5700 810.7150 999.5000 811.2850 ;
      RECT 900.5000 810.7150 920.0000 811.2850 ;
      RECT 99.8350 810.7150 119.5000 811.2850 ;
      RECT 20.5000 810.7150 99.2650 811.2850 ;
      RECT 900.5000 809.4850 999.5000 810.7150 ;
      RECT 20.5000 809.4850 119.5000 810.7150 ;
      RECT 920.5700 808.9150 999.5000 809.4850 ;
      RECT 900.5000 808.9150 920.0000 809.4850 ;
      RECT 99.8350 808.9150 119.5000 809.4850 ;
      RECT 20.5000 808.9150 99.2650 809.4850 ;
      RECT 900.5000 807.6850 999.5000 808.9150 ;
      RECT 20.5000 807.6850 119.5000 808.9150 ;
      RECT 920.5700 807.1150 999.5000 807.6850 ;
      RECT 900.5000 807.1150 920.0000 807.6850 ;
      RECT 99.8350 807.1150 119.5000 807.6850 ;
      RECT 20.5000 807.1150 99.2650 807.6850 ;
      RECT 900.5000 805.8850 999.5000 807.1150 ;
      RECT 20.5000 805.8850 119.5000 807.1150 ;
      RECT 920.5700 805.3150 999.5000 805.8850 ;
      RECT 900.5000 805.3150 920.0000 805.8850 ;
      RECT 99.8350 805.3150 119.5000 805.8850 ;
      RECT 20.5000 805.3150 99.2650 805.8850 ;
      RECT 900.5000 804.0850 999.5000 805.3150 ;
      RECT 20.5000 804.0850 119.5000 805.3150 ;
      RECT 920.5700 803.5150 999.5000 804.0850 ;
      RECT 900.5000 803.5150 920.0000 804.0850 ;
      RECT 99.8350 803.5150 119.5000 804.0850 ;
      RECT 20.5000 803.5150 99.2650 804.0850 ;
      RECT 900.5000 802.2850 999.5000 803.5150 ;
      RECT 20.5000 802.2850 119.5000 803.5150 ;
      RECT 920.5700 801.7150 999.5000 802.2850 ;
      RECT 900.5000 801.7150 920.0000 802.2850 ;
      RECT 99.8350 801.7150 119.5000 802.2850 ;
      RECT 20.5000 801.7150 99.2650 802.2850 ;
      RECT 900.5000 800.4850 999.5000 801.7150 ;
      RECT 20.5000 800.4850 119.5000 801.7150 ;
      RECT 920.5700 799.9150 999.5000 800.4850 ;
      RECT 900.5000 799.9150 920.0000 800.4850 ;
      RECT 99.8350 799.9150 119.5000 800.4850 ;
      RECT 20.5000 799.9150 99.2650 800.4850 ;
      RECT 900.5000 798.6850 999.5000 799.9150 ;
      RECT 20.5000 798.6850 119.5000 799.9150 ;
      RECT 920.5700 798.1150 999.5000 798.6850 ;
      RECT 900.5000 798.1150 920.0000 798.6850 ;
      RECT 99.8350 798.1150 119.5000 798.6850 ;
      RECT 20.5000 798.1150 99.2650 798.6850 ;
      RECT 900.5000 796.8850 999.5000 798.1150 ;
      RECT 20.5000 796.8850 119.5000 798.1150 ;
      RECT 920.5700 796.3150 999.5000 796.8850 ;
      RECT 900.5000 796.3150 920.0000 796.8850 ;
      RECT 99.8350 796.3150 119.5000 796.8850 ;
      RECT 20.5000 796.3150 99.2650 796.8850 ;
      RECT 900.5000 795.0850 999.5000 796.3150 ;
      RECT 20.5000 795.0850 119.5000 796.3150 ;
      RECT 920.5700 794.5150 999.5000 795.0850 ;
      RECT 900.5000 794.5150 920.0000 795.0850 ;
      RECT 99.8350 794.5150 119.5000 795.0850 ;
      RECT 20.5000 794.5150 99.2650 795.0850 ;
      RECT 900.5000 793.2850 999.5000 794.5150 ;
      RECT 20.5000 793.2850 119.5000 794.5150 ;
      RECT 920.5700 792.7150 999.5000 793.2850 ;
      RECT 900.5000 792.7150 920.0000 793.2850 ;
      RECT 99.8350 792.7150 119.5000 793.2850 ;
      RECT 20.5000 792.7150 99.2650 793.2850 ;
      RECT 900.5000 791.4850 999.5000 792.7150 ;
      RECT 20.5000 791.4850 119.5000 792.7150 ;
      RECT 920.5700 790.9150 999.5000 791.4850 ;
      RECT 900.5000 790.9150 920.0000 791.4850 ;
      RECT 99.8350 790.9150 119.5000 791.4850 ;
      RECT 20.5000 790.9150 99.2650 791.4850 ;
      RECT 900.5000 789.6850 999.5000 790.9150 ;
      RECT 20.5000 789.6850 119.5000 790.9150 ;
      RECT 920.5700 789.1150 999.5000 789.6850 ;
      RECT 900.5000 789.1150 920.0000 789.6850 ;
      RECT 99.8350 789.1150 119.5000 789.6850 ;
      RECT 20.5000 789.1150 99.2650 789.6850 ;
      RECT 900.5000 787.8850 999.5000 789.1150 ;
      RECT 20.5000 787.8850 119.5000 789.1150 ;
      RECT 920.5700 787.3150 999.5000 787.8850 ;
      RECT 900.5000 787.3150 920.0000 787.8850 ;
      RECT 99.8350 787.3150 119.5000 787.8850 ;
      RECT 20.5000 787.3150 99.2650 787.8850 ;
      RECT 900.5000 786.0850 999.5000 787.3150 ;
      RECT 20.5000 786.0850 119.5000 787.3150 ;
      RECT 920.5700 785.5150 999.5000 786.0850 ;
      RECT 900.5000 785.5150 920.0000 786.0850 ;
      RECT 99.8350 785.5150 119.5000 786.0850 ;
      RECT 20.5000 785.5150 99.2650 786.0850 ;
      RECT 900.5000 784.2850 999.5000 785.5150 ;
      RECT 20.5000 784.2850 119.5000 785.5150 ;
      RECT 920.5700 783.7150 999.5000 784.2850 ;
      RECT 900.5000 783.7150 920.0000 784.2850 ;
      RECT 99.8350 783.7150 119.5000 784.2850 ;
      RECT 20.5000 783.7150 99.2650 784.2850 ;
      RECT 900.5000 782.4850 999.5000 783.7150 ;
      RECT 20.5000 782.4850 119.5000 783.7150 ;
      RECT 920.5700 781.9150 999.5000 782.4850 ;
      RECT 900.5000 781.9150 920.0000 782.4850 ;
      RECT 99.8350 781.9150 119.5000 782.4850 ;
      RECT 20.5000 781.9150 99.2650 782.4850 ;
      RECT 900.5000 780.6850 999.5000 781.9150 ;
      RECT 20.5000 780.6850 119.5000 781.9150 ;
      RECT 920.5700 780.1150 999.5000 780.6850 ;
      RECT 900.5000 780.1150 920.0000 780.6850 ;
      RECT 99.8350 780.1150 119.5000 780.6850 ;
      RECT 20.5000 780.1150 99.2650 780.6850 ;
      RECT 900.5000 778.8850 999.5000 780.1150 ;
      RECT 20.5000 778.8850 119.5000 780.1150 ;
      RECT 920.5700 778.3150 999.5000 778.8850 ;
      RECT 900.5000 778.3150 920.0000 778.8850 ;
      RECT 99.8350 778.3150 119.5000 778.8850 ;
      RECT 20.5000 778.3150 99.2650 778.8850 ;
      RECT 900.5000 777.0850 999.5000 778.3150 ;
      RECT 20.5000 777.0850 119.5000 778.3150 ;
      RECT 920.5700 776.5150 999.5000 777.0850 ;
      RECT 900.5000 776.5150 920.0000 777.0850 ;
      RECT 99.8350 776.5150 119.5000 777.0850 ;
      RECT 20.5000 776.5150 99.2650 777.0850 ;
      RECT 900.5000 775.2850 999.5000 776.5150 ;
      RECT 20.5000 775.2850 119.5000 776.5150 ;
      RECT 920.5700 774.7150 999.5000 775.2850 ;
      RECT 900.5000 774.7150 920.0000 775.2850 ;
      RECT 99.8350 774.7150 119.5000 775.2850 ;
      RECT 20.5000 774.7150 99.2650 775.2850 ;
      RECT 900.5000 773.4850 999.5000 774.7150 ;
      RECT 20.5000 773.4850 119.5000 774.7150 ;
      RECT 920.5700 772.9150 999.5000 773.4850 ;
      RECT 900.5000 772.9150 920.0000 773.4850 ;
      RECT 99.8350 772.9150 119.5000 773.4850 ;
      RECT 20.5000 772.9150 99.2650 773.4850 ;
      RECT 900.5000 771.6850 999.5000 772.9150 ;
      RECT 20.5000 771.6850 119.5000 772.9150 ;
      RECT 920.5700 771.1150 999.5000 771.6850 ;
      RECT 900.5000 771.1150 920.0000 771.6850 ;
      RECT 99.8350 771.1150 119.5000 771.6850 ;
      RECT 20.5000 771.1150 99.2650 771.6850 ;
      RECT 900.5000 769.8850 999.5000 771.1150 ;
      RECT 20.5000 769.8850 119.5000 771.1150 ;
      RECT 920.5700 769.3150 999.5000 769.8850 ;
      RECT 900.5000 769.3150 920.0000 769.8850 ;
      RECT 99.8350 769.3150 119.5000 769.8850 ;
      RECT 20.5000 769.3150 99.2650 769.8850 ;
      RECT 900.5000 768.0850 999.5000 769.3150 ;
      RECT 20.5000 768.0850 119.5000 769.3150 ;
      RECT 920.5700 767.5150 999.5000 768.0850 ;
      RECT 900.5000 767.5150 920.0000 768.0850 ;
      RECT 99.8350 767.5150 119.5000 768.0850 ;
      RECT 20.5000 767.5150 99.2650 768.0850 ;
      RECT 900.5000 766.2850 999.5000 767.5150 ;
      RECT 20.5000 766.2850 119.5000 767.5150 ;
      RECT 920.5700 765.7150 999.5000 766.2850 ;
      RECT 900.5000 765.7150 920.0000 766.2850 ;
      RECT 99.8350 765.7150 119.5000 766.2850 ;
      RECT 20.5000 765.7150 99.2650 766.2850 ;
      RECT 900.5000 764.4850 999.5000 765.7150 ;
      RECT 20.5000 764.4850 119.5000 765.7150 ;
      RECT 920.5700 763.9150 999.5000 764.4850 ;
      RECT 900.5000 763.9150 920.0000 764.4850 ;
      RECT 99.8350 763.9150 119.5000 764.4850 ;
      RECT 20.5000 763.9150 99.2650 764.4850 ;
      RECT 900.5000 762.6850 999.5000 763.9150 ;
      RECT 20.5000 762.6850 119.5000 763.9150 ;
      RECT 920.5700 762.1150 999.5000 762.6850 ;
      RECT 900.5000 762.1150 920.0000 762.6850 ;
      RECT 99.8350 762.1150 119.5000 762.6850 ;
      RECT 20.5000 762.1150 99.2650 762.6850 ;
      RECT 900.5000 760.8850 999.5000 762.1150 ;
      RECT 20.5000 760.8850 119.5000 762.1150 ;
      RECT 920.5700 760.3150 999.5000 760.8850 ;
      RECT 900.5000 760.3150 920.0000 760.8850 ;
      RECT 99.8350 760.3150 119.5000 760.8850 ;
      RECT 20.5000 760.3150 99.2650 760.8850 ;
      RECT 900.5000 759.0850 999.5000 760.3150 ;
      RECT 20.5000 759.0850 119.5000 760.3150 ;
      RECT 920.5700 758.5150 999.5000 759.0850 ;
      RECT 900.5000 758.5150 920.0000 759.0850 ;
      RECT 99.8350 758.5150 119.5000 759.0850 ;
      RECT 20.5000 758.5150 99.2650 759.0850 ;
      RECT 900.5000 757.2850 999.5000 758.5150 ;
      RECT 20.5000 757.2850 119.5000 758.5150 ;
      RECT 920.5700 756.7150 999.5000 757.2850 ;
      RECT 900.5000 756.7150 920.0000 757.2850 ;
      RECT 99.8350 756.7150 119.5000 757.2850 ;
      RECT 20.5000 756.7150 99.2650 757.2850 ;
      RECT 900.5000 755.4850 999.5000 756.7150 ;
      RECT 20.5000 755.4850 119.5000 756.7150 ;
      RECT 920.5700 754.9150 999.5000 755.4850 ;
      RECT 900.5000 754.9150 920.0000 755.4850 ;
      RECT 99.8350 754.9150 119.5000 755.4850 ;
      RECT 20.5000 754.9150 99.2650 755.4850 ;
      RECT 900.5000 753.6850 999.5000 754.9150 ;
      RECT 20.5000 753.6850 119.5000 754.9150 ;
      RECT 920.5700 753.1150 999.5000 753.6850 ;
      RECT 900.5000 753.1150 920.0000 753.6850 ;
      RECT 99.8350 753.1150 119.5000 753.6850 ;
      RECT 20.5000 753.1150 99.2650 753.6850 ;
      RECT 900.5000 751.8850 999.5000 753.1150 ;
      RECT 20.5000 751.8850 119.5000 753.1150 ;
      RECT 920.5700 751.3150 999.5000 751.8850 ;
      RECT 900.5000 751.3150 920.0000 751.8850 ;
      RECT 99.8350 751.3150 119.5000 751.8850 ;
      RECT 20.5000 751.3150 99.2650 751.8850 ;
      RECT 900.5000 750.0850 999.5000 751.3150 ;
      RECT 20.5000 750.0850 119.5000 751.3150 ;
      RECT 920.5700 749.5150 999.5000 750.0850 ;
      RECT 900.5000 749.5150 920.0000 750.0850 ;
      RECT 99.8350 749.5150 119.5000 750.0850 ;
      RECT 20.5000 749.5150 99.2650 750.0850 ;
      RECT 900.5000 748.2850 999.5000 749.5150 ;
      RECT 20.5000 748.2850 119.5000 749.5150 ;
      RECT 920.5700 747.7150 999.5000 748.2850 ;
      RECT 900.5000 747.7150 920.0000 748.2850 ;
      RECT 99.8350 747.7150 119.5000 748.2850 ;
      RECT 20.5000 747.7150 99.2650 748.2850 ;
      RECT 900.5000 746.4850 999.5000 747.7150 ;
      RECT 20.5000 746.4850 119.5000 747.7150 ;
      RECT 920.5700 745.9150 999.5000 746.4850 ;
      RECT 900.5000 745.9150 920.0000 746.4850 ;
      RECT 99.8350 745.9150 119.5000 746.4850 ;
      RECT 20.5000 745.9150 99.2650 746.4850 ;
      RECT 900.5000 744.6850 999.5000 745.9150 ;
      RECT 20.5000 744.6850 119.5000 745.9150 ;
      RECT 920.5700 744.1150 999.5000 744.6850 ;
      RECT 900.5000 744.1150 920.0000 744.6850 ;
      RECT 99.8350 744.1150 119.5000 744.6850 ;
      RECT 20.5000 744.1150 99.2650 744.6850 ;
      RECT 900.5000 742.8850 999.5000 744.1150 ;
      RECT 20.5000 742.8850 119.5000 744.1150 ;
      RECT 920.5700 742.3150 999.5000 742.8850 ;
      RECT 900.5000 742.3150 920.0000 742.8850 ;
      RECT 99.8350 742.3150 119.5000 742.8850 ;
      RECT 20.5000 742.3150 99.2650 742.8850 ;
      RECT 900.5000 741.0850 999.5000 742.3150 ;
      RECT 20.5000 741.0850 119.5000 742.3150 ;
      RECT 920.5700 740.5150 999.5000 741.0850 ;
      RECT 900.5000 740.5150 920.0000 741.0850 ;
      RECT 99.8350 740.5150 119.5000 741.0850 ;
      RECT 20.5000 740.5150 99.2650 741.0850 ;
      RECT 900.5000 739.2850 999.5000 740.5150 ;
      RECT 20.5000 739.2850 119.5000 740.5150 ;
      RECT 920.5700 738.7150 999.5000 739.2850 ;
      RECT 900.5000 738.7150 920.0000 739.2850 ;
      RECT 99.8350 738.7150 119.5000 739.2850 ;
      RECT 20.5000 738.7150 99.2650 739.2850 ;
      RECT 900.5000 737.4850 999.5000 738.7150 ;
      RECT 20.5000 737.4850 119.5000 738.7150 ;
      RECT 920.5700 736.9150 999.5000 737.4850 ;
      RECT 900.5000 736.9150 920.0000 737.4850 ;
      RECT 99.8350 736.9150 119.5000 737.4850 ;
      RECT 20.5000 736.9150 99.2650 737.4850 ;
      RECT 900.5000 735.6850 999.5000 736.9150 ;
      RECT 20.5000 735.6850 119.5000 736.9150 ;
      RECT 920.5700 735.1150 999.5000 735.6850 ;
      RECT 900.5000 735.1150 920.0000 735.6850 ;
      RECT 99.8350 735.1150 119.5000 735.6850 ;
      RECT 20.5000 735.1150 99.2650 735.6850 ;
      RECT 900.5000 733.8850 999.5000 735.1150 ;
      RECT 20.5000 733.8850 119.5000 735.1150 ;
      RECT 920.5700 733.3150 999.5000 733.8850 ;
      RECT 900.5000 733.3150 920.0000 733.8850 ;
      RECT 99.8350 733.3150 119.5000 733.8850 ;
      RECT 20.5000 733.3150 99.2650 733.8850 ;
      RECT 900.5000 732.0850 999.5000 733.3150 ;
      RECT 20.5000 732.0850 119.5000 733.3150 ;
      RECT 920.5700 731.5150 999.5000 732.0850 ;
      RECT 900.5000 731.5150 920.0000 732.0850 ;
      RECT 99.8350 731.5150 119.5000 732.0850 ;
      RECT 20.5000 731.5150 99.2650 732.0850 ;
      RECT 900.5000 730.2850 999.5000 731.5150 ;
      RECT 20.5000 730.2850 119.5000 731.5150 ;
      RECT 920.5700 729.7150 999.5000 730.2850 ;
      RECT 900.5000 729.7150 920.0000 730.2850 ;
      RECT 99.8350 729.7150 119.5000 730.2850 ;
      RECT 20.5000 729.7150 99.2650 730.2850 ;
      RECT 900.5000 728.4850 999.5000 729.7150 ;
      RECT 20.5000 728.4850 119.5000 729.7150 ;
      RECT 920.5700 727.9150 999.5000 728.4850 ;
      RECT 900.5000 727.9150 920.0000 728.4850 ;
      RECT 99.8350 727.9150 119.5000 728.4850 ;
      RECT 20.5000 727.9150 99.2650 728.4850 ;
      RECT 900.5000 726.6850 999.5000 727.9150 ;
      RECT 20.5000 726.6850 119.5000 727.9150 ;
      RECT 920.5700 726.1150 999.5000 726.6850 ;
      RECT 900.5000 726.1150 920.0000 726.6850 ;
      RECT 99.8350 726.1150 119.5000 726.6850 ;
      RECT 20.5000 726.1150 99.2650 726.6850 ;
      RECT 900.5000 724.8850 999.5000 726.1150 ;
      RECT 20.5000 724.8850 119.5000 726.1150 ;
      RECT 920.5700 724.3150 999.5000 724.8850 ;
      RECT 900.5000 724.3150 920.0000 724.8850 ;
      RECT 99.8350 724.3150 119.5000 724.8850 ;
      RECT 20.5000 724.3150 99.2650 724.8850 ;
      RECT 900.5000 723.0850 999.5000 724.3150 ;
      RECT 20.5000 723.0850 119.5000 724.3150 ;
      RECT 920.5700 722.5150 999.5000 723.0850 ;
      RECT 900.5000 722.5150 920.0000 723.0850 ;
      RECT 99.8350 722.5150 119.5000 723.0850 ;
      RECT 20.5000 722.5150 99.2650 723.0850 ;
      RECT 900.5000 721.2850 999.5000 722.5150 ;
      RECT 20.5000 721.2850 119.5000 722.5150 ;
      RECT 920.5700 720.7150 999.5000 721.2850 ;
      RECT 900.5000 720.7150 920.0000 721.2850 ;
      RECT 99.8350 720.7150 119.5000 721.2850 ;
      RECT 20.5000 720.7150 99.2650 721.2850 ;
      RECT 900.5000 719.4850 999.5000 720.7150 ;
      RECT 20.5000 719.4850 119.5000 720.7150 ;
      RECT 920.5700 718.9150 999.5000 719.4850 ;
      RECT 900.5000 718.9150 920.0000 719.4850 ;
      RECT 99.8350 718.9150 119.5000 719.4850 ;
      RECT 20.5000 718.9150 99.2650 719.4850 ;
      RECT 900.5000 717.6850 999.5000 718.9150 ;
      RECT 20.5000 717.6850 119.5000 718.9150 ;
      RECT 920.5700 717.1150 999.5000 717.6850 ;
      RECT 900.5000 717.1150 920.0000 717.6850 ;
      RECT 99.8350 717.1150 119.5000 717.6850 ;
      RECT 20.5000 717.1150 99.2650 717.6850 ;
      RECT 900.5000 715.8850 999.5000 717.1150 ;
      RECT 20.5000 715.8850 119.5000 717.1150 ;
      RECT 920.5700 715.3150 999.5000 715.8850 ;
      RECT 900.5000 715.3150 920.0000 715.8850 ;
      RECT 99.8350 715.3150 119.5000 715.8850 ;
      RECT 20.5000 715.3150 99.2650 715.8850 ;
      RECT 900.5000 714.0850 999.5000 715.3150 ;
      RECT 20.5000 714.0850 119.5000 715.3150 ;
      RECT 920.5700 713.5150 999.5000 714.0850 ;
      RECT 900.5000 713.5150 920.0000 714.0850 ;
      RECT 99.8350 713.5150 119.5000 714.0850 ;
      RECT 20.5000 713.5150 99.2650 714.0850 ;
      RECT 900.5000 712.2850 999.5000 713.5150 ;
      RECT 20.5000 712.2850 119.5000 713.5150 ;
      RECT 920.5700 711.7150 999.5000 712.2850 ;
      RECT 900.5000 711.7150 920.0000 712.2850 ;
      RECT 99.8350 711.7150 119.5000 712.2850 ;
      RECT 20.5000 711.7150 99.2650 712.2850 ;
      RECT 900.5000 710.4850 999.5000 711.7150 ;
      RECT 20.5000 710.4850 119.5000 711.7150 ;
      RECT 920.5700 709.9150 999.5000 710.4850 ;
      RECT 900.5000 709.9150 920.0000 710.4850 ;
      RECT 99.8350 709.9150 119.5000 710.4850 ;
      RECT 20.5000 709.9150 99.2650 710.4850 ;
      RECT 900.5000 708.6850 999.5000 709.9150 ;
      RECT 20.5000 708.6850 119.5000 709.9150 ;
      RECT 920.5700 708.1150 999.5000 708.6850 ;
      RECT 900.5000 708.1150 920.0000 708.6850 ;
      RECT 99.8350 708.1150 119.5000 708.6850 ;
      RECT 20.5000 708.1150 99.2650 708.6850 ;
      RECT 900.5000 706.8850 999.5000 708.1150 ;
      RECT 20.5000 706.8850 119.5000 708.1150 ;
      RECT 920.5700 706.3150 999.5000 706.8850 ;
      RECT 900.5000 706.3150 920.0000 706.8850 ;
      RECT 99.8350 706.3150 119.5000 706.8850 ;
      RECT 20.5000 706.3150 99.2650 706.8850 ;
      RECT 900.5000 705.0850 999.5000 706.3150 ;
      RECT 20.5000 705.0850 119.5000 706.3150 ;
      RECT 920.5700 704.5150 999.5000 705.0850 ;
      RECT 900.5000 704.5150 920.0000 705.0850 ;
      RECT 99.8350 704.5150 119.5000 705.0850 ;
      RECT 20.5000 704.5150 99.2650 705.0850 ;
      RECT 900.5000 703.2850 999.5000 704.5150 ;
      RECT 20.5000 703.2850 119.5000 704.5150 ;
      RECT 920.5700 702.7150 999.5000 703.2850 ;
      RECT 900.5000 702.7150 920.0000 703.2850 ;
      RECT 99.8350 702.7150 119.5000 703.2850 ;
      RECT 20.5000 702.7150 99.2650 703.2850 ;
      RECT 900.5000 701.4850 999.5000 702.7150 ;
      RECT 20.5000 701.4850 119.5000 702.7150 ;
      RECT 920.5700 700.9150 999.5000 701.4850 ;
      RECT 900.5000 700.9150 920.0000 701.4850 ;
      RECT 99.8350 700.9150 119.5000 701.4850 ;
      RECT 20.5000 700.9150 99.2650 701.4850 ;
      RECT 900.5000 699.6850 999.5000 700.9150 ;
      RECT 20.5000 699.6850 119.5000 700.9150 ;
      RECT 920.5700 699.1150 999.5000 699.6850 ;
      RECT 900.5000 699.1150 920.0000 699.6850 ;
      RECT 99.8350 699.1150 119.5000 699.6850 ;
      RECT 20.5000 699.1150 99.2650 699.6850 ;
      RECT 900.5000 697.8850 999.5000 699.1150 ;
      RECT 20.5000 697.8850 119.5000 699.1150 ;
      RECT 920.5700 697.3150 999.5000 697.8850 ;
      RECT 900.5000 697.3150 920.0000 697.8850 ;
      RECT 99.8350 697.3150 119.5000 697.8850 ;
      RECT 20.5000 697.3150 99.2650 697.8850 ;
      RECT 900.5000 696.0850 999.5000 697.3150 ;
      RECT 20.5000 696.0850 119.5000 697.3150 ;
      RECT 920.5700 695.5150 999.5000 696.0850 ;
      RECT 900.5000 695.5150 920.0000 696.0850 ;
      RECT 99.8350 695.5150 119.5000 696.0850 ;
      RECT 20.5000 695.5150 99.2650 696.0850 ;
      RECT 900.5000 694.2850 999.5000 695.5150 ;
      RECT 20.5000 694.2850 119.5000 695.5150 ;
      RECT 920.5700 693.7150 999.5000 694.2850 ;
      RECT 900.5000 693.7150 920.0000 694.2850 ;
      RECT 99.8350 693.7150 119.5000 694.2850 ;
      RECT 20.5000 693.7150 99.2650 694.2850 ;
      RECT 900.5000 692.4850 999.5000 693.7150 ;
      RECT 20.5000 692.4850 119.5000 693.7150 ;
      RECT 920.5700 691.9150 999.5000 692.4850 ;
      RECT 900.5000 691.9150 920.0000 692.4850 ;
      RECT 99.8350 691.9150 119.5000 692.4850 ;
      RECT 20.5000 691.9150 99.2650 692.4850 ;
      RECT 900.5000 690.6850 999.5000 691.9150 ;
      RECT 20.5000 690.6850 119.5000 691.9150 ;
      RECT 920.5700 690.1150 999.5000 690.6850 ;
      RECT 900.5000 690.1150 920.0000 690.6850 ;
      RECT 99.8350 690.1150 119.5000 690.6850 ;
      RECT 20.5000 690.1150 99.2650 690.6850 ;
      RECT 900.5000 688.8850 999.5000 690.1150 ;
      RECT 20.5000 688.8850 119.5000 690.1150 ;
      RECT 920.5700 688.3150 999.5000 688.8850 ;
      RECT 900.5000 688.3150 920.0000 688.8850 ;
      RECT 99.8350 688.3150 119.5000 688.8850 ;
      RECT 20.5000 688.3150 99.2650 688.8850 ;
      RECT 900.5000 687.0850 999.5000 688.3150 ;
      RECT 20.5000 687.0850 119.5000 688.3150 ;
      RECT 920.5700 686.5150 999.5000 687.0850 ;
      RECT 900.5000 686.5150 920.0000 687.0850 ;
      RECT 99.8350 686.5150 119.5000 687.0850 ;
      RECT 20.5000 686.5150 99.2650 687.0850 ;
      RECT 900.5000 685.2850 999.5000 686.5150 ;
      RECT 20.5000 685.2850 119.5000 686.5150 ;
      RECT 920.5700 684.7150 999.5000 685.2850 ;
      RECT 900.5000 684.7150 920.0000 685.2850 ;
      RECT 99.8350 684.7150 119.5000 685.2850 ;
      RECT 20.5000 684.7150 99.2650 685.2850 ;
      RECT 900.5000 683.4850 999.5000 684.7150 ;
      RECT 20.5000 683.4850 119.5000 684.7150 ;
      RECT 920.5700 682.9150 999.5000 683.4850 ;
      RECT 900.5000 682.9150 920.0000 683.4850 ;
      RECT 99.8350 682.9150 119.5000 683.4850 ;
      RECT 20.5000 682.9150 99.2650 683.4850 ;
      RECT 900.5000 681.6850 999.5000 682.9150 ;
      RECT 20.5000 681.6850 119.5000 682.9150 ;
      RECT 920.5700 681.1150 999.5000 681.6850 ;
      RECT 900.5000 681.1150 920.0000 681.6850 ;
      RECT 99.8350 681.1150 119.5000 681.6850 ;
      RECT 20.5000 681.1150 99.2650 681.6850 ;
      RECT 900.5000 679.8850 999.5000 681.1150 ;
      RECT 20.5000 679.8850 119.5000 681.1150 ;
      RECT 920.5700 679.3150 999.5000 679.8850 ;
      RECT 900.5000 679.3150 920.0000 679.8850 ;
      RECT 99.8350 679.3150 119.5000 679.8850 ;
      RECT 20.5000 679.3150 99.2650 679.8850 ;
      RECT 900.5000 678.0850 999.5000 679.3150 ;
      RECT 20.5000 678.0850 119.5000 679.3150 ;
      RECT 920.5700 677.5150 999.5000 678.0850 ;
      RECT 900.5000 677.5150 920.0000 678.0850 ;
      RECT 99.8350 677.5150 119.5000 678.0850 ;
      RECT 20.5000 677.5150 99.2650 678.0850 ;
      RECT 900.5000 676.2850 999.5000 677.5150 ;
      RECT 20.5000 676.2850 119.5000 677.5150 ;
      RECT 920.5700 675.7150 999.5000 676.2850 ;
      RECT 900.5000 675.7150 920.0000 676.2850 ;
      RECT 99.8350 675.7150 119.5000 676.2850 ;
      RECT 20.5000 675.7150 99.2650 676.2850 ;
      RECT 900.5000 674.4850 999.5000 675.7150 ;
      RECT 20.5000 674.4850 119.5000 675.7150 ;
      RECT 920.5700 673.9150 999.5000 674.4850 ;
      RECT 900.5000 673.9150 920.0000 674.4850 ;
      RECT 99.8350 673.9150 119.5000 674.4850 ;
      RECT 20.5000 673.9150 99.2650 674.4850 ;
      RECT 900.5000 672.6850 999.5000 673.9150 ;
      RECT 20.5000 672.6850 119.5000 673.9150 ;
      RECT 920.5700 672.1150 999.5000 672.6850 ;
      RECT 900.5000 672.1150 920.0000 672.6850 ;
      RECT 99.8350 672.1150 119.5000 672.6850 ;
      RECT 20.5000 672.1150 99.2650 672.6850 ;
      RECT 900.5000 670.8850 999.5000 672.1150 ;
      RECT 20.5000 670.8850 119.5000 672.1150 ;
      RECT 920.5700 670.3150 999.5000 670.8850 ;
      RECT 900.5000 670.3150 920.0000 670.8850 ;
      RECT 99.8350 670.3150 119.5000 670.8850 ;
      RECT 20.5000 670.3150 99.2650 670.8850 ;
      RECT 900.5000 669.0850 999.5000 670.3150 ;
      RECT 20.5000 669.0850 119.5000 670.3150 ;
      RECT 920.5700 668.5150 999.5000 669.0850 ;
      RECT 900.5000 668.5150 920.0000 669.0850 ;
      RECT 99.8350 668.5150 119.5000 669.0850 ;
      RECT 20.5000 668.5150 99.2650 669.0850 ;
      RECT 900.5000 667.2850 999.5000 668.5150 ;
      RECT 20.5000 667.2850 119.5000 668.5150 ;
      RECT 920.5700 666.7150 999.5000 667.2850 ;
      RECT 900.5000 666.7150 920.0000 667.2850 ;
      RECT 99.8350 666.7150 119.5000 667.2850 ;
      RECT 20.5000 666.7150 99.2650 667.2850 ;
      RECT 900.5000 665.4850 999.5000 666.7150 ;
      RECT 20.5000 665.4850 119.5000 666.7150 ;
      RECT 920.5700 664.9150 999.5000 665.4850 ;
      RECT 900.5000 664.9150 920.0000 665.4850 ;
      RECT 99.8350 664.9150 119.5000 665.4850 ;
      RECT 20.5000 664.9150 99.2650 665.4850 ;
      RECT 900.5000 663.6850 999.5000 664.9150 ;
      RECT 20.5000 663.6850 119.5000 664.9150 ;
      RECT 920.5700 663.1150 999.5000 663.6850 ;
      RECT 900.5000 663.1150 920.0000 663.6850 ;
      RECT 99.8350 663.1150 119.5000 663.6850 ;
      RECT 20.5000 663.1150 99.2650 663.6850 ;
      RECT 900.5000 661.8850 999.5000 663.1150 ;
      RECT 20.5000 661.8850 119.5000 663.1150 ;
      RECT 920.5700 661.3150 999.5000 661.8850 ;
      RECT 900.5000 661.3150 920.0000 661.8850 ;
      RECT 99.8350 661.3150 119.5000 661.8850 ;
      RECT 20.5000 661.3150 99.2650 661.8850 ;
      RECT 900.5000 660.0850 999.5000 661.3150 ;
      RECT 20.5000 660.0850 119.5000 661.3150 ;
      RECT 920.5700 659.5150 999.5000 660.0850 ;
      RECT 900.5000 659.5150 920.0000 660.0850 ;
      RECT 99.8350 659.5150 119.5000 660.0850 ;
      RECT 20.5000 659.5150 99.2650 660.0850 ;
      RECT 900.5000 658.2850 999.5000 659.5150 ;
      RECT 20.5000 658.2850 119.5000 659.5150 ;
      RECT 920.5700 657.7150 999.5000 658.2850 ;
      RECT 900.5000 657.7150 920.0000 658.2850 ;
      RECT 99.8350 657.7150 119.5000 658.2850 ;
      RECT 20.5000 657.7150 99.2650 658.2850 ;
      RECT 900.5000 656.4850 999.5000 657.7150 ;
      RECT 20.5000 656.4850 119.5000 657.7150 ;
      RECT 920.5700 655.9150 999.5000 656.4850 ;
      RECT 900.5000 655.9150 920.0000 656.4850 ;
      RECT 99.8350 655.9150 119.5000 656.4850 ;
      RECT 20.5000 655.9150 99.2650 656.4850 ;
      RECT 900.5000 654.6850 999.5000 655.9150 ;
      RECT 20.5000 654.6850 119.5000 655.9150 ;
      RECT 920.5700 654.1150 999.5000 654.6850 ;
      RECT 900.5000 654.1150 920.0000 654.6850 ;
      RECT 99.8350 654.1150 119.5000 654.6850 ;
      RECT 20.5000 654.1150 99.2650 654.6850 ;
      RECT 900.5000 652.8850 999.5000 654.1150 ;
      RECT 20.5000 652.8850 119.5000 654.1150 ;
      RECT 920.5700 652.3150 999.5000 652.8850 ;
      RECT 900.5000 652.3150 920.0000 652.8850 ;
      RECT 99.8350 652.3150 119.5000 652.8850 ;
      RECT 20.5000 652.3150 99.2650 652.8850 ;
      RECT 900.5000 651.0850 999.5000 652.3150 ;
      RECT 20.5000 651.0850 119.5000 652.3150 ;
      RECT 920.5700 650.5150 999.5000 651.0850 ;
      RECT 900.5000 650.5150 920.0000 651.0850 ;
      RECT 99.8350 650.5150 119.5000 651.0850 ;
      RECT 20.5000 650.5150 99.2650 651.0850 ;
      RECT 900.5000 649.2850 999.5000 650.5150 ;
      RECT 20.5000 649.2850 119.5000 650.5150 ;
      RECT 920.5700 648.7150 999.5000 649.2850 ;
      RECT 900.5000 648.7150 920.0000 649.2850 ;
      RECT 99.8350 648.7150 119.5000 649.2850 ;
      RECT 20.5000 648.7150 99.2650 649.2850 ;
      RECT 900.5000 647.4850 999.5000 648.7150 ;
      RECT 20.5000 647.4850 119.5000 648.7150 ;
      RECT 920.5700 646.9150 999.5000 647.4850 ;
      RECT 900.5000 646.9150 920.0000 647.4850 ;
      RECT 99.8350 646.9150 119.5000 647.4850 ;
      RECT 20.5000 646.9150 99.2650 647.4850 ;
      RECT 900.5000 645.6850 999.5000 646.9150 ;
      RECT 20.5000 645.6850 119.5000 646.9150 ;
      RECT 920.5700 645.1150 999.5000 645.6850 ;
      RECT 900.5000 645.1150 920.0000 645.6850 ;
      RECT 99.8350 645.1150 119.5000 645.6850 ;
      RECT 20.5000 645.1150 99.2650 645.6850 ;
      RECT 900.5000 643.8850 999.5000 645.1150 ;
      RECT 20.5000 643.8850 119.5000 645.1150 ;
      RECT 920.5700 643.3150 999.5000 643.8850 ;
      RECT 900.5000 643.3150 920.0000 643.8850 ;
      RECT 99.8350 643.3150 119.5000 643.8850 ;
      RECT 20.5000 643.3150 99.2650 643.8850 ;
      RECT 900.5000 642.0850 999.5000 643.3150 ;
      RECT 20.5000 642.0850 119.5000 643.3150 ;
      RECT 920.5700 641.5150 999.5000 642.0850 ;
      RECT 900.5000 641.5150 920.0000 642.0850 ;
      RECT 99.8350 641.5150 119.5000 642.0850 ;
      RECT 20.5000 641.5150 99.2650 642.0850 ;
      RECT 900.5000 640.2850 999.5000 641.5150 ;
      RECT 20.5000 640.2850 119.5000 641.5150 ;
      RECT 920.5700 639.7150 999.5000 640.2850 ;
      RECT 900.5000 639.7150 920.0000 640.2850 ;
      RECT 99.8350 639.7150 119.5000 640.2850 ;
      RECT 20.5000 639.7150 99.2650 640.2850 ;
      RECT 900.5000 638.4850 999.5000 639.7150 ;
      RECT 20.5000 638.4850 119.5000 639.7150 ;
      RECT 920.5700 637.9150 999.5000 638.4850 ;
      RECT 900.5000 637.9150 920.0000 638.4850 ;
      RECT 99.8350 637.9150 119.5000 638.4850 ;
      RECT 20.5000 637.9150 99.2650 638.4850 ;
      RECT 900.5000 636.6850 999.5000 637.9150 ;
      RECT 20.5000 636.6850 119.5000 637.9150 ;
      RECT 920.5700 636.1150 999.5000 636.6850 ;
      RECT 900.5000 636.1150 920.0000 636.6850 ;
      RECT 99.8350 636.1150 119.5000 636.6850 ;
      RECT 20.5000 636.1150 99.2650 636.6850 ;
      RECT 900.5000 634.8850 999.5000 636.1150 ;
      RECT 20.5000 634.8850 119.5000 636.1150 ;
      RECT 920.5700 634.3150 999.5000 634.8850 ;
      RECT 900.5000 634.3150 920.0000 634.8850 ;
      RECT 99.8350 634.3150 119.5000 634.8850 ;
      RECT 20.5000 634.3150 99.2650 634.8850 ;
      RECT 900.5000 633.0850 999.5000 634.3150 ;
      RECT 20.5000 633.0850 119.5000 634.3150 ;
      RECT 920.5700 632.5150 999.5000 633.0850 ;
      RECT 900.5000 632.5150 920.0000 633.0850 ;
      RECT 99.8350 632.5150 119.5000 633.0850 ;
      RECT 20.5000 632.5150 99.2650 633.0850 ;
      RECT 900.5000 631.2850 999.5000 632.5150 ;
      RECT 20.5000 631.2850 119.5000 632.5150 ;
      RECT 920.5700 630.7150 999.5000 631.2850 ;
      RECT 900.5000 630.7150 920.0000 631.2850 ;
      RECT 99.8350 630.7150 119.5000 631.2850 ;
      RECT 20.5000 630.7150 99.2650 631.2850 ;
      RECT 900.5000 629.4850 999.5000 630.7150 ;
      RECT 20.5000 629.4850 119.5000 630.7150 ;
      RECT 920.5700 628.9150 999.5000 629.4850 ;
      RECT 900.5000 628.9150 920.0000 629.4850 ;
      RECT 99.8350 628.9150 119.5000 629.4850 ;
      RECT 20.5000 628.9150 99.2650 629.4850 ;
      RECT 900.5000 627.6850 999.5000 628.9150 ;
      RECT 20.5000 627.6850 119.5000 628.9150 ;
      RECT 920.5700 627.1150 999.5000 627.6850 ;
      RECT 900.5000 627.1150 920.0000 627.6850 ;
      RECT 99.8350 627.1150 119.5000 627.6850 ;
      RECT 20.5000 627.1150 99.2650 627.6850 ;
      RECT 900.5000 625.8850 999.5000 627.1150 ;
      RECT 20.5000 625.8850 119.5000 627.1150 ;
      RECT 920.5700 625.3150 999.5000 625.8850 ;
      RECT 900.5000 625.3150 920.0000 625.8850 ;
      RECT 99.8350 625.3150 119.5000 625.8850 ;
      RECT 20.5000 625.3150 99.2650 625.8850 ;
      RECT 900.5000 624.0850 999.5000 625.3150 ;
      RECT 20.5000 624.0850 119.5000 625.3150 ;
      RECT 920.5700 623.5150 999.5000 624.0850 ;
      RECT 900.5000 623.5150 920.0000 624.0850 ;
      RECT 99.8350 623.5150 119.5000 624.0850 ;
      RECT 20.5000 623.5150 99.2650 624.0850 ;
      RECT 900.5000 622.2850 999.5000 623.5150 ;
      RECT 20.5000 622.2850 119.5000 623.5150 ;
      RECT 920.5700 621.7150 999.5000 622.2850 ;
      RECT 900.5000 621.7150 920.0000 622.2850 ;
      RECT 99.8350 621.7150 119.5000 622.2850 ;
      RECT 20.5000 621.7150 99.2650 622.2850 ;
      RECT 900.5000 620.4850 999.5000 621.7150 ;
      RECT 20.5000 620.4850 119.5000 621.7150 ;
      RECT 920.5700 619.9150 999.5000 620.4850 ;
      RECT 900.5000 619.9150 920.0000 620.4850 ;
      RECT 99.8350 619.9150 119.5000 620.4850 ;
      RECT 20.5000 619.9150 99.2650 620.4850 ;
      RECT 900.5000 618.6850 999.5000 619.9150 ;
      RECT 20.5000 618.6850 119.5000 619.9150 ;
      RECT 920.5700 618.1150 999.5000 618.6850 ;
      RECT 900.5000 618.1150 920.0000 618.6850 ;
      RECT 99.8350 618.1150 119.5000 618.6850 ;
      RECT 20.5000 618.1150 99.2650 618.6850 ;
      RECT 900.5000 616.8850 999.5000 618.1150 ;
      RECT 20.5000 616.8850 119.5000 618.1150 ;
      RECT 920.5700 616.3150 999.5000 616.8850 ;
      RECT 900.5000 616.3150 920.0000 616.8850 ;
      RECT 99.8350 616.3150 119.5000 616.8850 ;
      RECT 20.5000 616.3150 99.2650 616.8850 ;
      RECT 900.5000 615.0850 999.5000 616.3150 ;
      RECT 20.5000 615.0850 119.5000 616.3150 ;
      RECT 920.5700 614.5150 999.5000 615.0850 ;
      RECT 900.5000 614.5150 920.0000 615.0850 ;
      RECT 99.8350 614.5150 119.5000 615.0850 ;
      RECT 20.5000 614.5150 99.2650 615.0850 ;
      RECT 900.5000 613.2850 999.5000 614.5150 ;
      RECT 20.5000 613.2850 119.5000 614.5150 ;
      RECT 920.5700 612.7150 999.5000 613.2850 ;
      RECT 900.5000 612.7150 920.0000 613.2850 ;
      RECT 99.8350 612.7150 119.5000 613.2850 ;
      RECT 20.5000 612.7150 99.2650 613.2850 ;
      RECT 900.5000 611.4850 999.5000 612.7150 ;
      RECT 20.5000 611.4850 119.5000 612.7150 ;
      RECT 920.5700 610.9150 999.5000 611.4850 ;
      RECT 900.5000 610.9150 920.0000 611.4850 ;
      RECT 99.8350 610.9150 119.5000 611.4850 ;
      RECT 20.5000 610.9150 99.2650 611.4850 ;
      RECT 900.5000 609.6850 999.5000 610.9150 ;
      RECT 20.5000 609.6850 119.5000 610.9150 ;
      RECT 920.5700 609.1150 999.5000 609.6850 ;
      RECT 900.5000 609.1150 920.0000 609.6850 ;
      RECT 99.8350 609.1150 119.5000 609.6850 ;
      RECT 20.5000 609.1150 99.2650 609.6850 ;
      RECT 900.5000 607.8850 999.5000 609.1150 ;
      RECT 20.5000 607.8850 119.5000 609.1150 ;
      RECT 920.5700 607.3150 999.5000 607.8850 ;
      RECT 900.5000 607.3150 920.0000 607.8850 ;
      RECT 99.8350 607.3150 119.5000 607.8850 ;
      RECT 20.5000 607.3150 99.2650 607.8850 ;
      RECT 900.5000 606.0850 999.5000 607.3150 ;
      RECT 20.5000 606.0850 119.5000 607.3150 ;
      RECT 920.5700 605.5150 999.5000 606.0850 ;
      RECT 900.5000 605.5150 920.0000 606.0850 ;
      RECT 99.8350 605.5150 119.5000 606.0850 ;
      RECT 20.5000 605.5150 99.2650 606.0850 ;
      RECT 900.5000 604.2850 999.5000 605.5150 ;
      RECT 20.5000 604.2850 119.5000 605.5150 ;
      RECT 920.5700 603.7150 999.5000 604.2850 ;
      RECT 900.5000 603.7150 920.0000 604.2850 ;
      RECT 99.8350 603.7150 119.5000 604.2850 ;
      RECT 20.5000 603.7150 99.2650 604.2850 ;
      RECT 900.5000 602.4850 999.5000 603.7150 ;
      RECT 20.5000 602.4850 119.5000 603.7150 ;
      RECT 920.5700 601.9150 999.5000 602.4850 ;
      RECT 900.5000 601.9150 920.0000 602.4850 ;
      RECT 99.8350 601.9150 119.5000 602.4850 ;
      RECT 20.5000 601.9150 99.2650 602.4850 ;
      RECT 900.5000 600.6850 999.5000 601.9150 ;
      RECT 20.5000 600.6850 119.5000 601.9150 ;
      RECT 920.5700 600.1150 999.5000 600.6850 ;
      RECT 900.5000 600.1150 920.0000 600.6850 ;
      RECT 99.8350 600.1150 119.5000 600.6850 ;
      RECT 20.5000 600.1150 99.2650 600.6850 ;
      RECT 900.5000 519.6850 999.5000 600.1150 ;
      RECT 20.5000 519.6850 119.5000 600.1150 ;
      RECT 920.5700 519.1150 999.5000 519.6850 ;
      RECT 900.5000 519.1150 920.0000 519.6850 ;
      RECT 99.8350 519.1150 119.5000 519.6850 ;
      RECT 20.5000 519.1150 99.2650 519.6850 ;
      RECT 900.5000 517.8850 999.5000 519.1150 ;
      RECT 20.5000 517.8850 119.5000 519.1150 ;
      RECT 920.5700 517.3150 999.5000 517.8850 ;
      RECT 900.5000 517.3150 920.0000 517.8850 ;
      RECT 99.8350 517.3150 119.5000 517.8850 ;
      RECT 20.5000 517.3150 99.2650 517.8850 ;
      RECT 900.5000 516.0850 999.5000 517.3150 ;
      RECT 20.5000 516.0850 119.5000 517.3150 ;
      RECT 920.5700 515.5150 999.5000 516.0850 ;
      RECT 900.5000 515.5150 920.0000 516.0850 ;
      RECT 99.8350 515.5150 119.5000 516.0850 ;
      RECT 20.5000 515.5150 99.2650 516.0850 ;
      RECT 900.5000 514.2850 999.5000 515.5150 ;
      RECT 20.5000 514.2850 119.5000 515.5150 ;
      RECT 920.5700 513.7150 999.5000 514.2850 ;
      RECT 900.5000 513.7150 920.0000 514.2850 ;
      RECT 99.8350 513.7150 119.5000 514.2850 ;
      RECT 20.5000 513.7150 99.2650 514.2850 ;
      RECT 900.5000 512.4850 999.5000 513.7150 ;
      RECT 20.5000 512.4850 119.5000 513.7150 ;
      RECT 920.5700 511.9150 999.5000 512.4850 ;
      RECT 900.5000 511.9150 920.0000 512.4850 ;
      RECT 99.8350 511.9150 119.5000 512.4850 ;
      RECT 20.5000 511.9150 99.2650 512.4850 ;
      RECT 900.5000 510.6850 999.5000 511.9150 ;
      RECT 20.5000 510.6850 119.5000 511.9150 ;
      RECT 920.5700 510.1150 999.5000 510.6850 ;
      RECT 900.5000 510.1150 920.0000 510.6850 ;
      RECT 99.8350 510.1150 119.5000 510.6850 ;
      RECT 20.5000 510.1150 99.2650 510.6850 ;
      RECT 900.5000 508.8850 999.5000 510.1150 ;
      RECT 20.5000 508.8850 119.5000 510.1150 ;
      RECT 920.5700 508.3150 999.5000 508.8850 ;
      RECT 900.5000 508.3150 920.0000 508.8850 ;
      RECT 99.8350 508.3150 119.5000 508.8850 ;
      RECT 20.5000 508.3150 99.2650 508.8850 ;
      RECT 900.5000 507.0850 999.5000 508.3150 ;
      RECT 20.5000 507.0850 119.5000 508.3150 ;
      RECT 920.5700 506.5150 999.5000 507.0850 ;
      RECT 900.5000 506.5150 920.0000 507.0850 ;
      RECT 99.8350 506.5150 119.5000 507.0850 ;
      RECT 20.5000 506.5150 99.2650 507.0850 ;
      RECT 900.5000 505.2850 999.5000 506.5150 ;
      RECT 20.5000 505.2850 119.5000 506.5150 ;
      RECT 920.5700 504.7150 999.5000 505.2850 ;
      RECT 900.5000 504.7150 920.0000 505.2850 ;
      RECT 99.8350 504.7150 119.5000 505.2850 ;
      RECT 20.5000 504.7150 99.2650 505.2850 ;
      RECT 900.5000 503.4850 999.5000 504.7150 ;
      RECT 20.5000 503.4850 119.5000 504.7150 ;
      RECT 920.5700 502.9150 999.5000 503.4850 ;
      RECT 900.5000 502.9150 920.0000 503.4850 ;
      RECT 99.8350 502.9150 119.5000 503.4850 ;
      RECT 20.5000 502.9150 99.2650 503.4850 ;
      RECT 900.5000 501.6850 999.5000 502.9150 ;
      RECT 20.5000 501.6850 119.5000 502.9150 ;
      RECT 920.5700 501.1150 999.5000 501.6850 ;
      RECT 900.5000 501.1150 920.0000 501.6850 ;
      RECT 99.8350 501.1150 119.5000 501.6850 ;
      RECT 20.5000 501.1150 99.2650 501.6850 ;
      RECT 900.5000 499.8850 999.5000 501.1150 ;
      RECT 20.5000 499.8850 119.5000 501.1150 ;
      RECT 920.5700 499.3150 999.5000 499.8850 ;
      RECT 900.5000 499.3150 920.0000 499.8850 ;
      RECT 99.8350 499.3150 119.5000 499.8850 ;
      RECT 20.5000 499.3150 99.2650 499.8850 ;
      RECT 900.5000 498.0850 999.5000 499.3150 ;
      RECT 20.5000 498.0850 119.5000 499.3150 ;
      RECT 920.5700 497.5150 999.5000 498.0850 ;
      RECT 900.5000 497.5150 920.0000 498.0850 ;
      RECT 99.8350 497.5150 119.5000 498.0850 ;
      RECT 20.5000 497.5150 99.2650 498.0850 ;
      RECT 900.5000 496.2850 999.5000 497.5150 ;
      RECT 20.5000 496.2850 119.5000 497.5150 ;
      RECT 920.5700 495.7150 999.5000 496.2850 ;
      RECT 900.5000 495.7150 920.0000 496.2850 ;
      RECT 99.8350 495.7150 119.5000 496.2850 ;
      RECT 20.5000 495.7150 99.2650 496.2850 ;
      RECT 900.5000 494.4850 999.5000 495.7150 ;
      RECT 20.5000 494.4850 119.5000 495.7150 ;
      RECT 920.5700 493.9150 999.5000 494.4850 ;
      RECT 900.5000 493.9150 920.0000 494.4850 ;
      RECT 99.8350 493.9150 119.5000 494.4850 ;
      RECT 20.5000 493.9150 99.2650 494.4850 ;
      RECT 900.5000 492.6850 999.5000 493.9150 ;
      RECT 20.5000 492.6850 119.5000 493.9150 ;
      RECT 920.5700 492.1150 999.5000 492.6850 ;
      RECT 900.5000 492.1150 920.0000 492.6850 ;
      RECT 99.8350 492.1150 119.5000 492.6850 ;
      RECT 20.5000 492.1150 99.2650 492.6850 ;
      RECT 900.5000 490.8850 999.5000 492.1150 ;
      RECT 20.5000 490.8850 119.5000 492.1150 ;
      RECT 920.5700 490.3150 999.5000 490.8850 ;
      RECT 900.5000 490.3150 920.0000 490.8850 ;
      RECT 99.8350 490.3150 119.5000 490.8850 ;
      RECT 20.5000 490.3150 99.2650 490.8850 ;
      RECT 900.5000 489.0850 999.5000 490.3150 ;
      RECT 20.5000 489.0850 119.5000 490.3150 ;
      RECT 920.5700 488.5150 999.5000 489.0850 ;
      RECT 900.5000 488.5150 920.0000 489.0850 ;
      RECT 99.8350 488.5150 119.5000 489.0850 ;
      RECT 20.5000 488.5150 99.2650 489.0850 ;
      RECT 900.5000 487.2850 999.5000 488.5150 ;
      RECT 20.5000 487.2850 119.5000 488.5150 ;
      RECT 920.5700 486.7150 999.5000 487.2850 ;
      RECT 900.5000 486.7150 920.0000 487.2850 ;
      RECT 99.8350 486.7150 119.5000 487.2850 ;
      RECT 20.5000 486.7150 99.2650 487.2850 ;
      RECT 900.5000 485.4850 999.5000 486.7150 ;
      RECT 20.5000 485.4850 119.5000 486.7150 ;
      RECT 920.5700 484.9150 999.5000 485.4850 ;
      RECT 900.5000 484.9150 920.0000 485.4850 ;
      RECT 99.8350 484.9150 119.5000 485.4850 ;
      RECT 20.5000 484.9150 99.2650 485.4850 ;
      RECT 900.5000 483.6850 999.5000 484.9150 ;
      RECT 20.5000 483.6850 119.5000 484.9150 ;
      RECT 920.5700 483.1150 999.5000 483.6850 ;
      RECT 900.5000 483.1150 920.0000 483.6850 ;
      RECT 99.8350 483.1150 119.5000 483.6850 ;
      RECT 20.5000 483.1150 99.2650 483.6850 ;
      RECT 900.5000 481.8850 999.5000 483.1150 ;
      RECT 20.5000 481.8850 119.5000 483.1150 ;
      RECT 920.5700 481.3150 999.5000 481.8850 ;
      RECT 900.5000 481.3150 920.0000 481.8850 ;
      RECT 99.8350 481.3150 119.5000 481.8850 ;
      RECT 20.5000 481.3150 99.2650 481.8850 ;
      RECT 900.5000 480.0850 999.5000 481.3150 ;
      RECT 20.5000 480.0850 119.5000 481.3150 ;
      RECT 920.5700 479.5150 999.5000 480.0850 ;
      RECT 900.5000 479.5150 920.0000 480.0850 ;
      RECT 99.8350 479.5150 119.5000 480.0850 ;
      RECT 20.5000 479.5150 99.2650 480.0850 ;
      RECT 900.5000 478.2850 999.5000 479.5150 ;
      RECT 20.5000 478.2850 119.5000 479.5150 ;
      RECT 920.5700 477.7150 999.5000 478.2850 ;
      RECT 900.5000 477.7150 920.0000 478.2850 ;
      RECT 99.8350 477.7150 119.5000 478.2850 ;
      RECT 20.5000 477.7150 99.2650 478.2850 ;
      RECT 900.5000 476.4850 999.5000 477.7150 ;
      RECT 20.5000 476.4850 119.5000 477.7150 ;
      RECT 920.5700 475.9150 999.5000 476.4850 ;
      RECT 900.5000 475.9150 920.0000 476.4850 ;
      RECT 99.8350 475.9150 119.5000 476.4850 ;
      RECT 20.5000 475.9150 99.2650 476.4850 ;
      RECT 900.5000 474.6850 999.5000 475.9150 ;
      RECT 20.5000 474.6850 119.5000 475.9150 ;
      RECT 920.5700 474.1150 999.5000 474.6850 ;
      RECT 900.5000 474.1150 920.0000 474.6850 ;
      RECT 99.8350 474.1150 119.5000 474.6850 ;
      RECT 20.5000 474.1150 99.2650 474.6850 ;
      RECT 900.5000 472.8850 999.5000 474.1150 ;
      RECT 20.5000 472.8850 119.5000 474.1150 ;
      RECT 920.5700 472.3150 999.5000 472.8850 ;
      RECT 900.5000 472.3150 920.0000 472.8850 ;
      RECT 99.8350 472.3150 119.5000 472.8850 ;
      RECT 20.5000 472.3150 99.2650 472.8850 ;
      RECT 900.5000 471.0850 999.5000 472.3150 ;
      RECT 20.5000 471.0850 119.5000 472.3150 ;
      RECT 920.5700 470.5150 999.5000 471.0850 ;
      RECT 900.5000 470.5150 920.0000 471.0850 ;
      RECT 99.8350 470.5150 119.5000 471.0850 ;
      RECT 20.5000 470.5150 99.2650 471.0850 ;
      RECT 900.5000 469.2850 999.5000 470.5150 ;
      RECT 20.5000 469.2850 119.5000 470.5150 ;
      RECT 920.5700 468.7150 999.5000 469.2850 ;
      RECT 900.5000 468.7150 920.0000 469.2850 ;
      RECT 99.8350 468.7150 119.5000 469.2850 ;
      RECT 20.5000 468.7150 99.2650 469.2850 ;
      RECT 900.5000 467.4850 999.5000 468.7150 ;
      RECT 20.5000 467.4850 119.5000 468.7150 ;
      RECT 920.5700 466.9150 999.5000 467.4850 ;
      RECT 900.5000 466.9150 920.0000 467.4850 ;
      RECT 99.8350 466.9150 119.5000 467.4850 ;
      RECT 20.5000 466.9150 99.2650 467.4850 ;
      RECT 900.5000 465.6850 999.5000 466.9150 ;
      RECT 20.5000 465.6850 119.5000 466.9150 ;
      RECT 920.5700 465.1150 999.5000 465.6850 ;
      RECT 900.5000 465.1150 920.0000 465.6850 ;
      RECT 99.8350 465.1150 119.5000 465.6850 ;
      RECT 20.5000 465.1150 99.2650 465.6850 ;
      RECT 900.5000 463.8850 999.5000 465.1150 ;
      RECT 20.5000 463.8850 119.5000 465.1150 ;
      RECT 920.5700 463.3150 999.5000 463.8850 ;
      RECT 900.5000 463.3150 920.0000 463.8850 ;
      RECT 99.8350 463.3150 119.5000 463.8850 ;
      RECT 20.5000 463.3150 99.2650 463.8850 ;
      RECT 900.5000 462.0850 999.5000 463.3150 ;
      RECT 20.5000 462.0850 119.5000 463.3150 ;
      RECT 920.5700 461.5150 999.5000 462.0850 ;
      RECT 900.5000 461.5150 920.0000 462.0850 ;
      RECT 99.8350 461.5150 119.5000 462.0850 ;
      RECT 20.5000 461.5150 99.2650 462.0850 ;
      RECT 900.5000 460.2850 999.5000 461.5150 ;
      RECT 20.5000 460.2850 119.5000 461.5150 ;
      RECT 920.5700 459.7150 999.5000 460.2850 ;
      RECT 900.5000 459.7150 920.0000 460.2850 ;
      RECT 99.8350 459.7150 119.5000 460.2850 ;
      RECT 20.5000 459.7150 99.2650 460.2850 ;
      RECT 900.5000 458.4850 999.5000 459.7150 ;
      RECT 20.5000 458.4850 119.5000 459.7150 ;
      RECT 920.5700 457.9150 999.5000 458.4850 ;
      RECT 900.5000 457.9150 920.0000 458.4850 ;
      RECT 99.8350 457.9150 119.5000 458.4850 ;
      RECT 20.5000 457.9150 99.2650 458.4850 ;
      RECT 900.5000 456.6850 999.5000 457.9150 ;
      RECT 20.5000 456.6850 119.5000 457.9150 ;
      RECT 920.5700 456.1150 999.5000 456.6850 ;
      RECT 900.5000 456.1150 920.0000 456.6850 ;
      RECT 99.8350 456.1150 119.5000 456.6850 ;
      RECT 20.5000 456.1150 99.2650 456.6850 ;
      RECT 900.5000 454.8850 999.5000 456.1150 ;
      RECT 20.5000 454.8850 119.5000 456.1150 ;
      RECT 920.5700 454.3150 999.5000 454.8850 ;
      RECT 900.5000 454.3150 920.0000 454.8850 ;
      RECT 99.8350 454.3150 119.5000 454.8850 ;
      RECT 20.5000 454.3150 99.2650 454.8850 ;
      RECT 900.5000 453.0850 999.5000 454.3150 ;
      RECT 20.5000 453.0850 119.5000 454.3150 ;
      RECT 920.5700 452.5150 999.5000 453.0850 ;
      RECT 900.5000 452.5150 920.0000 453.0850 ;
      RECT 99.8350 452.5150 119.5000 453.0850 ;
      RECT 20.5000 452.5150 99.2650 453.0850 ;
      RECT 900.5000 451.2850 999.5000 452.5150 ;
      RECT 20.5000 451.2850 119.5000 452.5150 ;
      RECT 920.5700 450.7150 999.5000 451.2850 ;
      RECT 900.5000 450.7150 920.0000 451.2850 ;
      RECT 99.8350 450.7150 119.5000 451.2850 ;
      RECT 20.5000 450.7150 99.2650 451.2850 ;
      RECT 900.5000 449.4850 999.5000 450.7150 ;
      RECT 20.5000 449.4850 119.5000 450.7150 ;
      RECT 920.5700 448.9150 999.5000 449.4850 ;
      RECT 900.5000 448.9150 920.0000 449.4850 ;
      RECT 99.8350 448.9150 119.5000 449.4850 ;
      RECT 20.5000 448.9150 99.2650 449.4850 ;
      RECT 900.5000 447.6850 999.5000 448.9150 ;
      RECT 20.5000 447.6850 119.5000 448.9150 ;
      RECT 920.5700 447.1150 999.5000 447.6850 ;
      RECT 900.5000 447.1150 920.0000 447.6850 ;
      RECT 99.8350 447.1150 119.5000 447.6850 ;
      RECT 20.5000 447.1150 99.2650 447.6850 ;
      RECT 900.5000 445.8850 999.5000 447.1150 ;
      RECT 20.5000 445.8850 119.5000 447.1150 ;
      RECT 920.5700 445.3150 999.5000 445.8850 ;
      RECT 900.5000 445.3150 920.0000 445.8850 ;
      RECT 99.8350 445.3150 119.5000 445.8850 ;
      RECT 20.5000 445.3150 99.2650 445.8850 ;
      RECT 900.5000 444.0850 999.5000 445.3150 ;
      RECT 20.5000 444.0850 119.5000 445.3150 ;
      RECT 920.5700 443.5150 999.5000 444.0850 ;
      RECT 900.5000 443.5150 920.0000 444.0850 ;
      RECT 99.8350 443.5150 119.5000 444.0850 ;
      RECT 20.5000 443.5150 99.2650 444.0850 ;
      RECT 900.5000 442.2850 999.5000 443.5150 ;
      RECT 20.5000 442.2850 119.5000 443.5150 ;
      RECT 920.5700 441.7150 999.5000 442.2850 ;
      RECT 900.5000 441.7150 920.0000 442.2850 ;
      RECT 99.8350 441.7150 119.5000 442.2850 ;
      RECT 20.5000 441.7150 99.2650 442.2850 ;
      RECT 900.5000 440.4850 999.5000 441.7150 ;
      RECT 20.5000 440.4850 119.5000 441.7150 ;
      RECT 920.5700 439.9150 999.5000 440.4850 ;
      RECT 900.5000 439.9150 920.0000 440.4850 ;
      RECT 99.8350 439.9150 119.5000 440.4850 ;
      RECT 20.5000 439.9150 99.2650 440.4850 ;
      RECT 900.5000 438.6850 999.5000 439.9150 ;
      RECT 20.5000 438.6850 119.5000 439.9150 ;
      RECT 920.5700 438.1150 999.5000 438.6850 ;
      RECT 900.5000 438.1150 920.0000 438.6850 ;
      RECT 99.8350 438.1150 119.5000 438.6850 ;
      RECT 20.5000 438.1150 99.2650 438.6850 ;
      RECT 900.5000 436.8850 999.5000 438.1150 ;
      RECT 20.5000 436.8850 119.5000 438.1150 ;
      RECT 920.5700 436.3150 999.5000 436.8850 ;
      RECT 900.5000 436.3150 920.0000 436.8850 ;
      RECT 99.8350 436.3150 119.5000 436.8850 ;
      RECT 20.5000 436.3150 99.2650 436.8850 ;
      RECT 900.5000 435.0850 999.5000 436.3150 ;
      RECT 20.5000 435.0850 119.5000 436.3150 ;
      RECT 920.5700 434.5150 999.5000 435.0850 ;
      RECT 900.5000 434.5150 920.0000 435.0850 ;
      RECT 99.8350 434.5150 119.5000 435.0850 ;
      RECT 20.5000 434.5150 99.2650 435.0850 ;
      RECT 900.5000 433.2850 999.5000 434.5150 ;
      RECT 20.5000 433.2850 119.5000 434.5150 ;
      RECT 920.5700 432.7150 999.5000 433.2850 ;
      RECT 900.5000 432.7150 920.0000 433.2850 ;
      RECT 99.8350 432.7150 119.5000 433.2850 ;
      RECT 20.5000 432.7150 99.2650 433.2850 ;
      RECT 900.5000 431.4850 999.5000 432.7150 ;
      RECT 20.5000 431.4850 119.5000 432.7150 ;
      RECT 920.5700 430.9150 999.5000 431.4850 ;
      RECT 900.5000 430.9150 920.0000 431.4850 ;
      RECT 99.8350 430.9150 119.5000 431.4850 ;
      RECT 20.5000 430.9150 99.2650 431.4850 ;
      RECT 900.5000 429.6850 999.5000 430.9150 ;
      RECT 20.5000 429.6850 119.5000 430.9150 ;
      RECT 920.5700 429.1150 999.5000 429.6850 ;
      RECT 900.5000 429.1150 920.0000 429.6850 ;
      RECT 99.8350 429.1150 119.5000 429.6850 ;
      RECT 20.5000 429.1150 99.2650 429.6850 ;
      RECT 900.5000 427.8850 999.5000 429.1150 ;
      RECT 20.5000 427.8850 119.5000 429.1150 ;
      RECT 920.5700 427.3150 999.5000 427.8850 ;
      RECT 900.5000 427.3150 920.0000 427.8850 ;
      RECT 99.8350 427.3150 119.5000 427.8850 ;
      RECT 20.5000 427.3150 99.2650 427.8850 ;
      RECT 900.5000 426.0850 999.5000 427.3150 ;
      RECT 20.5000 426.0850 119.5000 427.3150 ;
      RECT 920.5700 425.5150 999.5000 426.0850 ;
      RECT 900.5000 425.5150 920.0000 426.0850 ;
      RECT 99.8350 425.5150 119.5000 426.0850 ;
      RECT 20.5000 425.5150 99.2650 426.0850 ;
      RECT 900.5000 424.2850 999.5000 425.5150 ;
      RECT 20.5000 424.2850 119.5000 425.5150 ;
      RECT 920.5700 423.7150 999.5000 424.2850 ;
      RECT 900.5000 423.7150 920.0000 424.2850 ;
      RECT 99.8350 423.7150 119.5000 424.2850 ;
      RECT 20.5000 423.7150 99.2650 424.2850 ;
      RECT 900.5000 422.4850 999.5000 423.7150 ;
      RECT 20.5000 422.4850 119.5000 423.7150 ;
      RECT 920.5700 421.9150 999.5000 422.4850 ;
      RECT 900.5000 421.9150 920.0000 422.4850 ;
      RECT 99.8350 421.9150 119.5000 422.4850 ;
      RECT 20.5000 421.9150 99.2650 422.4850 ;
      RECT 900.5000 420.6850 999.5000 421.9150 ;
      RECT 20.5000 420.6850 119.5000 421.9150 ;
      RECT 920.5700 420.1150 999.5000 420.6850 ;
      RECT 900.5000 420.1150 920.0000 420.6850 ;
      RECT 99.8350 420.1150 119.5000 420.6850 ;
      RECT 20.5000 420.1150 99.2650 420.6850 ;
      RECT 900.5000 418.8850 999.5000 420.1150 ;
      RECT 20.5000 418.8850 119.5000 420.1150 ;
      RECT 920.5700 418.3150 999.5000 418.8850 ;
      RECT 900.5000 418.3150 920.0000 418.8850 ;
      RECT 99.8350 418.3150 119.5000 418.8850 ;
      RECT 20.5000 418.3150 99.2650 418.8850 ;
      RECT 900.5000 417.0850 999.5000 418.3150 ;
      RECT 20.5000 417.0850 119.5000 418.3150 ;
      RECT 920.5700 416.5150 999.5000 417.0850 ;
      RECT 900.5000 416.5150 920.0000 417.0850 ;
      RECT 99.8350 416.5150 119.5000 417.0850 ;
      RECT 20.5000 416.5150 99.2650 417.0850 ;
      RECT 900.5000 415.2850 999.5000 416.5150 ;
      RECT 20.5000 415.2850 119.5000 416.5150 ;
      RECT 920.5700 414.7150 999.5000 415.2850 ;
      RECT 900.5000 414.7150 920.0000 415.2850 ;
      RECT 99.8350 414.7150 119.5000 415.2850 ;
      RECT 20.5000 414.7150 99.2650 415.2850 ;
      RECT 900.5000 413.4850 999.5000 414.7150 ;
      RECT 20.5000 413.4850 119.5000 414.7150 ;
      RECT 920.5700 412.9150 999.5000 413.4850 ;
      RECT 900.5000 412.9150 920.0000 413.4850 ;
      RECT 99.8350 412.9150 119.5000 413.4850 ;
      RECT 20.5000 412.9150 99.2650 413.4850 ;
      RECT 900.5000 411.6850 999.5000 412.9150 ;
      RECT 20.5000 411.6850 119.5000 412.9150 ;
      RECT 920.5700 411.1150 999.5000 411.6850 ;
      RECT 900.5000 411.1150 920.0000 411.6850 ;
      RECT 99.8350 411.1150 119.5000 411.6850 ;
      RECT 20.5000 411.1150 99.2650 411.6850 ;
      RECT 900.5000 409.8850 999.5000 411.1150 ;
      RECT 20.5000 409.8850 119.5000 411.1150 ;
      RECT 920.5700 409.3150 999.5000 409.8850 ;
      RECT 900.5000 409.3150 920.0000 409.8850 ;
      RECT 99.8350 409.3150 119.5000 409.8850 ;
      RECT 20.5000 409.3150 99.2650 409.8850 ;
      RECT 900.5000 408.0850 999.5000 409.3150 ;
      RECT 20.5000 408.0850 119.5000 409.3150 ;
      RECT 920.5700 407.5150 999.5000 408.0850 ;
      RECT 900.5000 407.5150 920.0000 408.0850 ;
      RECT 99.8350 407.5150 119.5000 408.0850 ;
      RECT 20.5000 407.5150 99.2650 408.0850 ;
      RECT 900.5000 406.2850 999.5000 407.5150 ;
      RECT 20.5000 406.2850 119.5000 407.5150 ;
      RECT 920.5700 405.7150 999.5000 406.2850 ;
      RECT 900.5000 405.7150 920.0000 406.2850 ;
      RECT 99.8350 405.7150 119.5000 406.2850 ;
      RECT 20.5000 405.7150 99.2650 406.2850 ;
      RECT 900.5000 404.4850 999.5000 405.7150 ;
      RECT 20.5000 404.4850 119.5000 405.7150 ;
      RECT 920.5700 403.9150 999.5000 404.4850 ;
      RECT 900.5000 403.9150 920.0000 404.4850 ;
      RECT 99.8350 403.9150 119.5000 404.4850 ;
      RECT 20.5000 403.9150 99.2650 404.4850 ;
      RECT 900.5000 402.6850 999.5000 403.9150 ;
      RECT 20.5000 402.6850 119.5000 403.9150 ;
      RECT 920.5700 402.1150 999.5000 402.6850 ;
      RECT 900.5000 402.1150 920.0000 402.6850 ;
      RECT 99.8350 402.1150 119.5000 402.6850 ;
      RECT 20.5000 402.1150 99.2650 402.6850 ;
      RECT 900.5000 400.8850 999.5000 402.1150 ;
      RECT 20.5000 400.8850 119.5000 402.1150 ;
      RECT 920.5700 400.3150 999.5000 400.8850 ;
      RECT 900.5000 400.3150 920.0000 400.8850 ;
      RECT 99.8350 400.3150 119.5000 400.8850 ;
      RECT 20.5000 400.3150 99.2650 400.8850 ;
      RECT 900.5000 399.0850 999.5000 400.3150 ;
      RECT 20.5000 399.0850 119.5000 400.3150 ;
      RECT 920.5700 398.5150 999.5000 399.0850 ;
      RECT 900.5000 398.5150 920.0000 399.0850 ;
      RECT 99.8350 398.5150 119.5000 399.0850 ;
      RECT 20.5000 398.5150 99.2650 399.0850 ;
      RECT 900.5000 397.2850 999.5000 398.5150 ;
      RECT 20.5000 397.2850 119.5000 398.5150 ;
      RECT 920.5700 396.7150 999.5000 397.2850 ;
      RECT 900.5000 396.7150 920.0000 397.2850 ;
      RECT 99.8350 396.7150 119.5000 397.2850 ;
      RECT 20.5000 396.7150 99.2650 397.2850 ;
      RECT 900.5000 395.4850 999.5000 396.7150 ;
      RECT 20.5000 395.4850 119.5000 396.7150 ;
      RECT 920.5700 394.9150 999.5000 395.4850 ;
      RECT 900.5000 394.9150 920.0000 395.4850 ;
      RECT 99.8350 394.9150 119.5000 395.4850 ;
      RECT 20.5000 394.9150 99.2650 395.4850 ;
      RECT 900.5000 393.6850 999.5000 394.9150 ;
      RECT 20.5000 393.6850 119.5000 394.9150 ;
      RECT 920.5700 393.1150 999.5000 393.6850 ;
      RECT 900.5000 393.1150 920.0000 393.6850 ;
      RECT 99.8350 393.1150 119.5000 393.6850 ;
      RECT 20.5000 393.1150 99.2650 393.6850 ;
      RECT 900.5000 391.8850 999.5000 393.1150 ;
      RECT 20.5000 391.8850 119.5000 393.1150 ;
      RECT 920.5700 391.3150 999.5000 391.8850 ;
      RECT 900.5000 391.3150 920.0000 391.8850 ;
      RECT 99.8350 391.3150 119.5000 391.8850 ;
      RECT 20.5000 391.3150 99.2650 391.8850 ;
      RECT 900.5000 390.0850 999.5000 391.3150 ;
      RECT 20.5000 390.0850 119.5000 391.3150 ;
      RECT 920.5700 389.5150 999.5000 390.0850 ;
      RECT 900.5000 389.5150 920.0000 390.0850 ;
      RECT 99.8350 389.5150 119.5000 390.0850 ;
      RECT 20.5000 389.5150 99.2650 390.0850 ;
      RECT 900.5000 388.2850 999.5000 389.5150 ;
      RECT 20.5000 388.2850 119.5000 389.5150 ;
      RECT 920.5700 387.7150 999.5000 388.2850 ;
      RECT 900.5000 387.7150 920.0000 388.2850 ;
      RECT 99.8350 387.7150 119.5000 388.2850 ;
      RECT 20.5000 387.7150 99.2650 388.2850 ;
      RECT 900.5000 386.4850 999.5000 387.7150 ;
      RECT 20.5000 386.4850 119.5000 387.7150 ;
      RECT 920.5700 385.9150 999.5000 386.4850 ;
      RECT 900.5000 385.9150 920.0000 386.4850 ;
      RECT 99.8350 385.9150 119.5000 386.4850 ;
      RECT 20.5000 385.9150 99.2650 386.4850 ;
      RECT 900.5000 384.6850 999.5000 385.9150 ;
      RECT 20.5000 384.6850 119.5000 385.9150 ;
      RECT 920.5700 384.1150 999.5000 384.6850 ;
      RECT 900.5000 384.1150 920.0000 384.6850 ;
      RECT 99.8350 384.1150 119.5000 384.6850 ;
      RECT 20.5000 384.1150 99.2650 384.6850 ;
      RECT 900.5000 382.8850 999.5000 384.1150 ;
      RECT 20.5000 382.8850 119.5000 384.1150 ;
      RECT 920.5700 382.3150 999.5000 382.8850 ;
      RECT 900.5000 382.3150 920.0000 382.8850 ;
      RECT 99.8350 382.3150 119.5000 382.8850 ;
      RECT 20.5000 382.3150 99.2650 382.8850 ;
      RECT 900.5000 381.0850 999.5000 382.3150 ;
      RECT 20.5000 381.0850 119.5000 382.3150 ;
      RECT 920.5700 380.5150 999.5000 381.0850 ;
      RECT 900.5000 380.5150 920.0000 381.0850 ;
      RECT 99.8350 380.5150 119.5000 381.0850 ;
      RECT 20.5000 380.5150 99.2650 381.0850 ;
      RECT 900.5000 379.2850 999.5000 380.5150 ;
      RECT 20.5000 379.2850 119.5000 380.5150 ;
      RECT 920.5700 378.7150 999.5000 379.2850 ;
      RECT 900.5000 378.7150 920.0000 379.2850 ;
      RECT 99.8350 378.7150 119.5000 379.2850 ;
      RECT 20.5000 378.7150 99.2650 379.2850 ;
      RECT 900.5000 377.4850 999.5000 378.7150 ;
      RECT 20.5000 377.4850 119.5000 378.7150 ;
      RECT 920.5700 376.9150 999.5000 377.4850 ;
      RECT 900.5000 376.9150 920.0000 377.4850 ;
      RECT 99.8350 376.9150 119.5000 377.4850 ;
      RECT 20.5000 376.9150 99.2650 377.4850 ;
      RECT 900.5000 375.6850 999.5000 376.9150 ;
      RECT 20.5000 375.6850 119.5000 376.9150 ;
      RECT 920.5700 375.1150 999.5000 375.6850 ;
      RECT 900.5000 375.1150 920.0000 375.6850 ;
      RECT 99.8350 375.1150 119.5000 375.6850 ;
      RECT 20.5000 375.1150 99.2650 375.6850 ;
      RECT 900.5000 373.8850 999.5000 375.1150 ;
      RECT 20.5000 373.8850 119.5000 375.1150 ;
      RECT 920.5700 373.3150 999.5000 373.8850 ;
      RECT 900.5000 373.3150 920.0000 373.8850 ;
      RECT 99.8350 373.3150 119.5000 373.8850 ;
      RECT 20.5000 373.3150 99.2650 373.8850 ;
      RECT 900.5000 372.0850 999.5000 373.3150 ;
      RECT 20.5000 372.0850 119.5000 373.3150 ;
      RECT 920.5700 371.5150 999.5000 372.0850 ;
      RECT 900.5000 371.5150 920.0000 372.0850 ;
      RECT 99.8350 371.5150 119.5000 372.0850 ;
      RECT 20.5000 371.5150 99.2650 372.0850 ;
      RECT 900.5000 370.2850 999.5000 371.5150 ;
      RECT 20.5000 370.2850 119.5000 371.5150 ;
      RECT 920.5700 369.7150 999.5000 370.2850 ;
      RECT 900.5000 369.7150 920.0000 370.2850 ;
      RECT 99.8350 369.7150 119.5000 370.2850 ;
      RECT 20.5000 369.7150 99.2650 370.2850 ;
      RECT 900.5000 368.4850 999.5000 369.7150 ;
      RECT 20.5000 368.4850 119.5000 369.7150 ;
      RECT 920.5700 367.9150 999.5000 368.4850 ;
      RECT 900.5000 367.9150 920.0000 368.4850 ;
      RECT 99.8350 367.9150 119.5000 368.4850 ;
      RECT 20.5000 367.9150 99.2650 368.4850 ;
      RECT 900.5000 366.6850 999.5000 367.9150 ;
      RECT 20.5000 366.6850 119.5000 367.9150 ;
      RECT 920.5700 366.1150 999.5000 366.6850 ;
      RECT 900.5000 366.1150 920.0000 366.6850 ;
      RECT 99.8350 366.1150 119.5000 366.6850 ;
      RECT 20.5000 366.1150 99.2650 366.6850 ;
      RECT 900.5000 364.8850 999.5000 366.1150 ;
      RECT 20.5000 364.8850 119.5000 366.1150 ;
      RECT 920.5700 364.3150 999.5000 364.8850 ;
      RECT 900.5000 364.3150 920.0000 364.8850 ;
      RECT 99.8350 364.3150 119.5000 364.8850 ;
      RECT 20.5000 364.3150 99.2650 364.8850 ;
      RECT 900.5000 363.0850 999.5000 364.3150 ;
      RECT 20.5000 363.0850 119.5000 364.3150 ;
      RECT 920.5700 362.5150 999.5000 363.0850 ;
      RECT 900.5000 362.5150 920.0000 363.0850 ;
      RECT 99.8350 362.5150 119.5000 363.0850 ;
      RECT 20.5000 362.5150 99.2650 363.0850 ;
      RECT 900.5000 361.2850 999.5000 362.5150 ;
      RECT 20.5000 361.2850 119.5000 362.5150 ;
      RECT 920.5700 360.7150 999.5000 361.2850 ;
      RECT 900.5000 360.7150 920.0000 361.2850 ;
      RECT 99.8350 360.7150 119.5000 361.2850 ;
      RECT 20.5000 360.7150 99.2650 361.2850 ;
      RECT 900.5000 359.4850 999.5000 360.7150 ;
      RECT 20.5000 359.4850 119.5000 360.7150 ;
      RECT 920.5700 358.9150 999.5000 359.4850 ;
      RECT 900.5000 358.9150 920.0000 359.4850 ;
      RECT 99.8350 358.9150 119.5000 359.4850 ;
      RECT 20.5000 358.9150 99.2650 359.4850 ;
      RECT 900.5000 357.6850 999.5000 358.9150 ;
      RECT 20.5000 357.6850 119.5000 358.9150 ;
      RECT 920.5700 357.1150 999.5000 357.6850 ;
      RECT 900.5000 357.1150 920.0000 357.6850 ;
      RECT 99.8350 357.1150 119.5000 357.6850 ;
      RECT 20.5000 357.1150 99.2650 357.6850 ;
      RECT 900.5000 355.8850 999.5000 357.1150 ;
      RECT 20.5000 355.8850 119.5000 357.1150 ;
      RECT 920.5700 355.3150 999.5000 355.8850 ;
      RECT 900.5000 355.3150 920.0000 355.8850 ;
      RECT 99.8350 355.3150 119.5000 355.8850 ;
      RECT 20.5000 355.3150 99.2650 355.8850 ;
      RECT 900.5000 354.0850 999.5000 355.3150 ;
      RECT 20.5000 354.0850 119.5000 355.3150 ;
      RECT 920.5700 353.5150 999.5000 354.0850 ;
      RECT 900.5000 353.5150 920.0000 354.0850 ;
      RECT 99.8350 353.5150 119.5000 354.0850 ;
      RECT 20.5000 353.5150 99.2650 354.0850 ;
      RECT 900.5000 352.2850 999.5000 353.5150 ;
      RECT 20.5000 352.2850 119.5000 353.5150 ;
      RECT 920.5700 351.7150 999.5000 352.2850 ;
      RECT 900.5000 351.7150 920.0000 352.2850 ;
      RECT 99.8350 351.7150 119.5000 352.2850 ;
      RECT 20.5000 351.7150 99.2650 352.2850 ;
      RECT 900.5000 350.4850 999.5000 351.7150 ;
      RECT 20.5000 350.4850 119.5000 351.7150 ;
      RECT 920.5700 349.9150 999.5000 350.4850 ;
      RECT 900.5000 349.9150 920.0000 350.4850 ;
      RECT 99.8350 349.9150 119.5000 350.4850 ;
      RECT 20.5000 349.9150 99.2650 350.4850 ;
      RECT 900.5000 348.6850 999.5000 349.9150 ;
      RECT 20.5000 348.6850 119.5000 349.9150 ;
      RECT 920.5700 348.1150 999.5000 348.6850 ;
      RECT 900.5000 348.1150 920.0000 348.6850 ;
      RECT 99.8350 348.1150 119.5000 348.6850 ;
      RECT 20.5000 348.1150 99.2650 348.6850 ;
      RECT 900.5000 346.8850 999.5000 348.1150 ;
      RECT 20.5000 346.8850 119.5000 348.1150 ;
      RECT 920.5700 346.3150 999.5000 346.8850 ;
      RECT 900.5000 346.3150 920.0000 346.8850 ;
      RECT 99.8350 346.3150 119.5000 346.8850 ;
      RECT 20.5000 346.3150 99.2650 346.8850 ;
      RECT 900.5000 345.0850 999.5000 346.3150 ;
      RECT 20.5000 345.0850 119.5000 346.3150 ;
      RECT 920.5700 344.5150 999.5000 345.0850 ;
      RECT 900.5000 344.5150 920.0000 345.0850 ;
      RECT 99.8350 344.5150 119.5000 345.0850 ;
      RECT 20.5000 344.5150 99.2650 345.0850 ;
      RECT 900.5000 343.2850 999.5000 344.5150 ;
      RECT 20.5000 343.2850 119.5000 344.5150 ;
      RECT 920.5700 342.7150 999.5000 343.2850 ;
      RECT 900.5000 342.7150 920.0000 343.2850 ;
      RECT 99.8350 342.7150 119.5000 343.2850 ;
      RECT 20.5000 342.7150 99.2650 343.2850 ;
      RECT 900.5000 341.4850 999.5000 342.7150 ;
      RECT 20.5000 341.4850 119.5000 342.7150 ;
      RECT 920.5700 340.9150 999.5000 341.4850 ;
      RECT 900.5000 340.9150 920.0000 341.4850 ;
      RECT 99.8350 340.9150 119.5000 341.4850 ;
      RECT 20.5000 340.9150 99.2650 341.4850 ;
      RECT 900.5000 339.6850 999.5000 340.9150 ;
      RECT 20.5000 339.6850 119.5000 340.9150 ;
      RECT 920.5700 339.1150 999.5000 339.6850 ;
      RECT 900.5000 339.1150 920.0000 339.6850 ;
      RECT 99.8350 339.1150 119.5000 339.6850 ;
      RECT 20.5000 339.1150 99.2650 339.6850 ;
      RECT 900.5000 337.8850 999.5000 339.1150 ;
      RECT 20.5000 337.8850 119.5000 339.1150 ;
      RECT 920.5700 337.3150 999.5000 337.8850 ;
      RECT 900.5000 337.3150 920.0000 337.8850 ;
      RECT 99.8350 337.3150 119.5000 337.8850 ;
      RECT 20.5000 337.3150 99.2650 337.8850 ;
      RECT 900.5000 336.0850 999.5000 337.3150 ;
      RECT 20.5000 336.0850 119.5000 337.3150 ;
      RECT 920.5700 335.5150 999.5000 336.0850 ;
      RECT 900.5000 335.5150 920.0000 336.0850 ;
      RECT 99.8350 335.5150 119.5000 336.0850 ;
      RECT 20.5000 335.5150 99.2650 336.0850 ;
      RECT 900.5000 334.2850 999.5000 335.5150 ;
      RECT 20.5000 334.2850 119.5000 335.5150 ;
      RECT 920.5700 333.7150 999.5000 334.2850 ;
      RECT 900.5000 333.7150 920.0000 334.2850 ;
      RECT 99.8350 333.7150 119.5000 334.2850 ;
      RECT 20.5000 333.7150 99.2650 334.2850 ;
      RECT 900.5000 332.4850 999.5000 333.7150 ;
      RECT 20.5000 332.4850 119.5000 333.7150 ;
      RECT 920.5700 331.9150 999.5000 332.4850 ;
      RECT 900.5000 331.9150 920.0000 332.4850 ;
      RECT 99.8350 331.9150 119.5000 332.4850 ;
      RECT 20.5000 331.9150 99.2650 332.4850 ;
      RECT 900.5000 330.6850 999.5000 331.9150 ;
      RECT 20.5000 330.6850 119.5000 331.9150 ;
      RECT 920.5700 330.1150 999.5000 330.6850 ;
      RECT 900.5000 330.1150 920.0000 330.6850 ;
      RECT 99.8350 330.1150 119.5000 330.6850 ;
      RECT 20.5000 330.1150 99.2650 330.6850 ;
      RECT 900.5000 328.8850 999.5000 330.1150 ;
      RECT 20.5000 328.8850 119.5000 330.1150 ;
      RECT 920.5700 328.3150 999.5000 328.8850 ;
      RECT 900.5000 328.3150 920.0000 328.8850 ;
      RECT 99.8350 328.3150 119.5000 328.8850 ;
      RECT 20.5000 328.3150 99.2650 328.8850 ;
      RECT 900.5000 327.0850 999.5000 328.3150 ;
      RECT 20.5000 327.0850 119.5000 328.3150 ;
      RECT 920.5700 326.5150 999.5000 327.0850 ;
      RECT 900.5000 326.5150 920.0000 327.0850 ;
      RECT 99.8350 326.5150 119.5000 327.0850 ;
      RECT 20.5000 326.5150 99.2650 327.0850 ;
      RECT 900.5000 325.2850 999.5000 326.5150 ;
      RECT 20.5000 325.2850 119.5000 326.5150 ;
      RECT 920.5700 324.7150 999.5000 325.2850 ;
      RECT 900.5000 324.7150 920.0000 325.2850 ;
      RECT 99.8350 324.7150 119.5000 325.2850 ;
      RECT 20.5000 324.7150 99.2650 325.2850 ;
      RECT 900.5000 323.4850 999.5000 324.7150 ;
      RECT 20.5000 323.4850 119.5000 324.7150 ;
      RECT 920.5700 322.9150 999.5000 323.4850 ;
      RECT 900.5000 322.9150 920.0000 323.4850 ;
      RECT 99.8350 322.9150 119.5000 323.4850 ;
      RECT 20.5000 322.9150 99.2650 323.4850 ;
      RECT 900.5000 321.6850 999.5000 322.9150 ;
      RECT 20.5000 321.6850 119.5000 322.9150 ;
      RECT 920.5700 321.1150 999.5000 321.6850 ;
      RECT 900.5000 321.1150 920.0000 321.6850 ;
      RECT 99.8350 321.1150 119.5000 321.6850 ;
      RECT 20.5000 321.1150 99.2650 321.6850 ;
      RECT 900.5000 319.8850 999.5000 321.1150 ;
      RECT 20.5000 319.8850 119.5000 321.1150 ;
      RECT 920.5700 319.3150 999.5000 319.8850 ;
      RECT 900.5000 319.3150 920.0000 319.8850 ;
      RECT 99.8350 319.3150 119.5000 319.8850 ;
      RECT 20.5000 319.3150 99.2650 319.8850 ;
      RECT 900.5000 318.0850 999.5000 319.3150 ;
      RECT 20.5000 318.0850 119.5000 319.3150 ;
      RECT 920.5700 317.5150 999.5000 318.0850 ;
      RECT 900.5000 317.5150 920.0000 318.0850 ;
      RECT 99.8350 317.5150 119.5000 318.0850 ;
      RECT 20.5000 317.5150 99.2650 318.0850 ;
      RECT 900.5000 316.2850 999.5000 317.5150 ;
      RECT 20.5000 316.2850 119.5000 317.5150 ;
      RECT 920.5700 315.7150 999.5000 316.2850 ;
      RECT 900.5000 315.7150 920.0000 316.2850 ;
      RECT 99.8350 315.7150 119.5000 316.2850 ;
      RECT 20.5000 315.7150 99.2650 316.2850 ;
      RECT 900.5000 314.4850 999.5000 315.7150 ;
      RECT 20.5000 314.4850 119.5000 315.7150 ;
      RECT 920.5700 313.9150 999.5000 314.4850 ;
      RECT 900.5000 313.9150 920.0000 314.4850 ;
      RECT 99.8350 313.9150 119.5000 314.4850 ;
      RECT 20.5000 313.9150 99.2650 314.4850 ;
      RECT 900.5000 312.6850 999.5000 313.9150 ;
      RECT 20.5000 312.6850 119.5000 313.9150 ;
      RECT 920.5700 312.1150 999.5000 312.6850 ;
      RECT 900.5000 312.1150 920.0000 312.6850 ;
      RECT 99.8350 312.1150 119.5000 312.6850 ;
      RECT 20.5000 312.1150 99.2650 312.6850 ;
      RECT 900.5000 310.8850 999.5000 312.1150 ;
      RECT 20.5000 310.8850 119.5000 312.1150 ;
      RECT 920.5700 310.3150 999.5000 310.8850 ;
      RECT 900.5000 310.3150 920.0000 310.8850 ;
      RECT 99.8350 310.3150 119.5000 310.8850 ;
      RECT 20.5000 310.3150 99.2650 310.8850 ;
      RECT 900.5000 309.0850 999.5000 310.3150 ;
      RECT 20.5000 309.0850 119.5000 310.3150 ;
      RECT 920.5700 308.5150 999.5000 309.0850 ;
      RECT 900.5000 308.5150 920.0000 309.0850 ;
      RECT 99.8350 308.5150 119.5000 309.0850 ;
      RECT 20.5000 308.5150 99.2650 309.0850 ;
      RECT 900.5000 307.2850 999.5000 308.5150 ;
      RECT 20.5000 307.2850 119.5000 308.5150 ;
      RECT 920.5700 306.7150 999.5000 307.2850 ;
      RECT 900.5000 306.7150 920.0000 307.2850 ;
      RECT 99.8350 306.7150 119.5000 307.2850 ;
      RECT 20.5000 306.7150 99.2650 307.2850 ;
      RECT 900.5000 305.4850 999.5000 306.7150 ;
      RECT 20.5000 305.4850 119.5000 306.7150 ;
      RECT 920.5700 304.9150 999.5000 305.4850 ;
      RECT 900.5000 304.9150 920.0000 305.4850 ;
      RECT 99.8350 304.9150 119.5000 305.4850 ;
      RECT 20.5000 304.9150 99.2650 305.4850 ;
      RECT 900.5000 303.6850 999.5000 304.9150 ;
      RECT 20.5000 303.6850 119.5000 304.9150 ;
      RECT 920.5700 303.1150 999.5000 303.6850 ;
      RECT 900.5000 303.1150 920.0000 303.6850 ;
      RECT 99.8350 303.1150 119.5000 303.6850 ;
      RECT 20.5000 303.1150 99.2650 303.6850 ;
      RECT 900.5000 301.8850 999.5000 303.1150 ;
      RECT 20.5000 301.8850 119.5000 303.1150 ;
      RECT 920.5700 301.3150 999.5000 301.8850 ;
      RECT 900.5000 301.3150 920.0000 301.8850 ;
      RECT 99.8350 301.3150 119.5000 301.8850 ;
      RECT 20.5000 301.3150 99.2650 301.8850 ;
      RECT 900.5000 300.0850 999.5000 301.3150 ;
      RECT 20.5000 300.0850 119.5000 301.3150 ;
      RECT 920.5700 299.5150 999.5000 300.0850 ;
      RECT 900.5000 299.5150 920.0000 300.0850 ;
      RECT 99.8350 299.5150 119.5000 300.0850 ;
      RECT 20.5000 299.5150 99.2650 300.0850 ;
      RECT 900.5000 298.2850 999.5000 299.5150 ;
      RECT 20.5000 298.2850 119.5000 299.5150 ;
      RECT 920.5700 297.7150 999.5000 298.2850 ;
      RECT 900.5000 297.7150 920.0000 298.2850 ;
      RECT 99.8350 297.7150 119.5000 298.2850 ;
      RECT 20.5000 297.7150 99.2650 298.2850 ;
      RECT 900.5000 296.4850 999.5000 297.7150 ;
      RECT 20.5000 296.4850 119.5000 297.7150 ;
      RECT 920.5700 295.9150 999.5000 296.4850 ;
      RECT 900.5000 295.9150 920.0000 296.4850 ;
      RECT 99.8350 295.9150 119.5000 296.4850 ;
      RECT 20.5000 295.9150 99.2650 296.4850 ;
      RECT 900.5000 294.6850 999.5000 295.9150 ;
      RECT 20.5000 294.6850 119.5000 295.9150 ;
      RECT 920.5700 294.1150 999.5000 294.6850 ;
      RECT 900.5000 294.1150 920.0000 294.6850 ;
      RECT 99.8350 294.1150 119.5000 294.6850 ;
      RECT 20.5000 294.1150 99.2650 294.6850 ;
      RECT 900.5000 292.8850 999.5000 294.1150 ;
      RECT 20.5000 292.8850 119.5000 294.1150 ;
      RECT 920.5700 292.3150 999.5000 292.8850 ;
      RECT 900.5000 292.3150 920.0000 292.8850 ;
      RECT 99.8350 292.3150 119.5000 292.8850 ;
      RECT 20.5000 292.3150 99.2650 292.8850 ;
      RECT 900.5000 291.0850 999.5000 292.3150 ;
      RECT 20.5000 291.0850 119.5000 292.3150 ;
      RECT 920.5700 290.5150 999.5000 291.0850 ;
      RECT 900.5000 290.5150 920.0000 291.0850 ;
      RECT 99.8350 290.5150 119.5000 291.0850 ;
      RECT 20.5000 290.5150 99.2650 291.0850 ;
      RECT 900.5000 289.2850 999.5000 290.5150 ;
      RECT 20.5000 289.2850 119.5000 290.5150 ;
      RECT 920.5700 288.7150 999.5000 289.2850 ;
      RECT 900.5000 288.7150 920.0000 289.2850 ;
      RECT 99.8350 288.7150 119.5000 289.2850 ;
      RECT 20.5000 288.7150 99.2650 289.2850 ;
      RECT 900.5000 287.4850 999.5000 288.7150 ;
      RECT 20.5000 287.4850 119.5000 288.7150 ;
      RECT 920.5700 286.9150 999.5000 287.4850 ;
      RECT 900.5000 286.9150 920.0000 287.4850 ;
      RECT 99.8350 286.9150 119.5000 287.4850 ;
      RECT 20.5000 286.9150 99.2650 287.4850 ;
      RECT 900.5000 285.6850 999.5000 286.9150 ;
      RECT 20.5000 285.6850 119.5000 286.9150 ;
      RECT 920.5700 285.1150 999.5000 285.6850 ;
      RECT 900.5000 285.1150 920.0000 285.6850 ;
      RECT 99.8350 285.1150 119.5000 285.6850 ;
      RECT 20.5000 285.1150 99.2650 285.6850 ;
      RECT 900.5000 283.8850 999.5000 285.1150 ;
      RECT 20.5000 283.8850 119.5000 285.1150 ;
      RECT 920.5700 283.3150 999.5000 283.8850 ;
      RECT 900.5000 283.3150 920.0000 283.8850 ;
      RECT 99.8350 283.3150 119.5000 283.8850 ;
      RECT 20.5000 283.3150 99.2650 283.8850 ;
      RECT 900.5000 282.0850 999.5000 283.3150 ;
      RECT 20.5000 282.0850 119.5000 283.3150 ;
      RECT 920.5700 281.5150 999.5000 282.0850 ;
      RECT 900.5000 281.5150 920.0000 282.0850 ;
      RECT 99.8350 281.5150 119.5000 282.0850 ;
      RECT 20.5000 281.5150 99.2650 282.0850 ;
      RECT 900.5000 280.2850 999.5000 281.5150 ;
      RECT 20.5000 280.2850 119.5000 281.5150 ;
      RECT 920.5700 279.7150 999.5000 280.2850 ;
      RECT 900.5000 279.7150 920.0000 280.2850 ;
      RECT 99.8350 279.7150 119.5000 280.2850 ;
      RECT 20.5000 279.7150 99.2650 280.2850 ;
      RECT 900.5000 278.4850 999.5000 279.7150 ;
      RECT 20.5000 278.4850 119.5000 279.7150 ;
      RECT 920.5700 277.9150 999.5000 278.4850 ;
      RECT 900.5000 277.9150 920.0000 278.4850 ;
      RECT 99.8350 277.9150 119.5000 278.4850 ;
      RECT 20.5000 277.9150 99.2650 278.4850 ;
      RECT 900.5000 276.6850 999.5000 277.9150 ;
      RECT 20.5000 276.6850 119.5000 277.9150 ;
      RECT 920.5700 276.1150 999.5000 276.6850 ;
      RECT 900.5000 276.1150 920.0000 276.6850 ;
      RECT 99.8350 276.1150 119.5000 276.6850 ;
      RECT 20.5000 276.1150 99.2650 276.6850 ;
      RECT 900.5000 274.8850 999.5000 276.1150 ;
      RECT 20.5000 274.8850 119.5000 276.1150 ;
      RECT 920.5700 274.3150 999.5000 274.8850 ;
      RECT 900.5000 274.3150 920.0000 274.8850 ;
      RECT 99.8350 274.3150 119.5000 274.8850 ;
      RECT 20.5000 274.3150 99.2650 274.8850 ;
      RECT 900.5000 273.0850 999.5000 274.3150 ;
      RECT 20.5000 273.0850 119.5000 274.3150 ;
      RECT 920.5700 272.5150 999.5000 273.0850 ;
      RECT 900.5000 272.5150 920.0000 273.0850 ;
      RECT 99.8350 272.5150 119.5000 273.0850 ;
      RECT 20.5000 272.5150 99.2650 273.0850 ;
      RECT 900.5000 271.2850 999.5000 272.5150 ;
      RECT 20.5000 271.2850 119.5000 272.5150 ;
      RECT 920.5700 270.7150 999.5000 271.2850 ;
      RECT 900.5000 270.7150 920.0000 271.2850 ;
      RECT 99.8350 270.7150 119.5000 271.2850 ;
      RECT 20.5000 270.7150 99.2650 271.2850 ;
      RECT 900.5000 269.4850 999.5000 270.7150 ;
      RECT 20.5000 269.4850 119.5000 270.7150 ;
      RECT 920.5700 268.9150 999.5000 269.4850 ;
      RECT 900.5000 268.9150 920.0000 269.4850 ;
      RECT 99.8350 268.9150 119.5000 269.4850 ;
      RECT 20.5000 268.9150 99.2650 269.4850 ;
      RECT 900.5000 267.6850 999.5000 268.9150 ;
      RECT 20.5000 267.6850 119.5000 268.9150 ;
      RECT 920.5700 267.1150 999.5000 267.6850 ;
      RECT 900.5000 267.1150 920.0000 267.6850 ;
      RECT 99.8350 267.1150 119.5000 267.6850 ;
      RECT 20.5000 267.1150 99.2650 267.6850 ;
      RECT 900.5000 265.8850 999.5000 267.1150 ;
      RECT 20.5000 265.8850 119.5000 267.1150 ;
      RECT 920.5700 265.3150 999.5000 265.8850 ;
      RECT 900.5000 265.3150 920.0000 265.8850 ;
      RECT 99.8350 265.3150 119.5000 265.8850 ;
      RECT 20.5000 265.3150 99.2650 265.8850 ;
      RECT 900.5000 264.0850 999.5000 265.3150 ;
      RECT 20.5000 264.0850 119.5000 265.3150 ;
      RECT 920.5700 263.5150 999.5000 264.0850 ;
      RECT 900.5000 263.5150 920.0000 264.0850 ;
      RECT 99.8350 263.5150 119.5000 264.0850 ;
      RECT 20.5000 263.5150 99.2650 264.0850 ;
      RECT 900.5000 262.2850 999.5000 263.5150 ;
      RECT 20.5000 262.2850 119.5000 263.5150 ;
      RECT 920.5700 261.7150 999.5000 262.2850 ;
      RECT 900.5000 261.7150 920.0000 262.2850 ;
      RECT 99.8350 261.7150 119.5000 262.2850 ;
      RECT 20.5000 261.7150 99.2650 262.2850 ;
      RECT 900.5000 260.4850 999.5000 261.7150 ;
      RECT 20.5000 260.4850 119.5000 261.7150 ;
      RECT 920.5700 259.9150 999.5000 260.4850 ;
      RECT 900.5000 259.9150 920.0000 260.4850 ;
      RECT 99.8350 259.9150 119.5000 260.4850 ;
      RECT 20.5000 259.9150 99.2650 260.4850 ;
      RECT 900.5000 258.6850 999.5000 259.9150 ;
      RECT 20.5000 258.6850 119.5000 259.9150 ;
      RECT 920.5700 258.1150 999.5000 258.6850 ;
      RECT 900.5000 258.1150 920.0000 258.6850 ;
      RECT 99.8350 258.1150 119.5000 258.6850 ;
      RECT 20.5000 258.1150 99.2650 258.6850 ;
      RECT 900.5000 256.8850 999.5000 258.1150 ;
      RECT 20.5000 256.8850 119.5000 258.1150 ;
      RECT 920.5700 256.3150 999.5000 256.8850 ;
      RECT 900.5000 256.3150 920.0000 256.8850 ;
      RECT 99.8350 256.3150 119.5000 256.8850 ;
      RECT 20.5000 256.3150 99.2650 256.8850 ;
      RECT 900.5000 255.0850 999.5000 256.3150 ;
      RECT 20.5000 255.0850 119.5000 256.3150 ;
      RECT 920.5700 254.5150 999.5000 255.0850 ;
      RECT 900.5000 254.5150 920.0000 255.0850 ;
      RECT 99.8350 254.5150 119.5000 255.0850 ;
      RECT 20.5000 254.5150 99.2650 255.0850 ;
      RECT 900.5000 253.2850 999.5000 254.5150 ;
      RECT 20.5000 253.2850 119.5000 254.5150 ;
      RECT 920.5700 252.7150 999.5000 253.2850 ;
      RECT 900.5000 252.7150 920.0000 253.2850 ;
      RECT 99.8350 252.7150 119.5000 253.2850 ;
      RECT 20.5000 252.7150 99.2650 253.2850 ;
      RECT 900.5000 251.4850 999.5000 252.7150 ;
      RECT 20.5000 251.4850 119.5000 252.7150 ;
      RECT 920.5700 250.9150 999.5000 251.4850 ;
      RECT 900.5000 250.9150 920.0000 251.4850 ;
      RECT 99.8350 250.9150 119.5000 251.4850 ;
      RECT 20.5000 250.9150 99.2650 251.4850 ;
      RECT 900.5000 249.6850 999.5000 250.9150 ;
      RECT 20.5000 249.6850 119.5000 250.9150 ;
      RECT 920.5700 249.1150 999.5000 249.6850 ;
      RECT 900.5000 249.1150 920.0000 249.6850 ;
      RECT 99.8350 249.1150 119.5000 249.6850 ;
      RECT 20.5000 249.1150 99.2650 249.6850 ;
      RECT 900.5000 247.8850 999.5000 249.1150 ;
      RECT 20.5000 247.8850 119.5000 249.1150 ;
      RECT 920.5700 247.3150 999.5000 247.8850 ;
      RECT 900.5000 247.3150 920.0000 247.8850 ;
      RECT 99.8350 247.3150 119.5000 247.8850 ;
      RECT 20.5000 247.3150 99.2650 247.8850 ;
      RECT 900.5000 246.0850 999.5000 247.3150 ;
      RECT 20.5000 246.0850 119.5000 247.3150 ;
      RECT 920.5700 245.5150 999.5000 246.0850 ;
      RECT 900.5000 245.5150 920.0000 246.0850 ;
      RECT 99.8350 245.5150 119.5000 246.0850 ;
      RECT 20.5000 245.5150 99.2650 246.0850 ;
      RECT 900.5000 244.2850 999.5000 245.5150 ;
      RECT 20.5000 244.2850 119.5000 245.5150 ;
      RECT 920.5700 243.7150 999.5000 244.2850 ;
      RECT 900.5000 243.7150 920.0000 244.2850 ;
      RECT 99.8350 243.7150 119.5000 244.2850 ;
      RECT 20.5000 243.7150 99.2650 244.2850 ;
      RECT 900.5000 242.4850 999.5000 243.7150 ;
      RECT 20.5000 242.4850 119.5000 243.7150 ;
      RECT 920.5700 241.9150 999.5000 242.4850 ;
      RECT 900.5000 241.9150 920.0000 242.4850 ;
      RECT 99.8350 241.9150 119.5000 242.4850 ;
      RECT 20.5000 241.9150 99.2650 242.4850 ;
      RECT 900.5000 240.6850 999.5000 241.9150 ;
      RECT 20.5000 240.6850 119.5000 241.9150 ;
      RECT 920.5700 240.1150 999.5000 240.6850 ;
      RECT 900.5000 240.1150 920.0000 240.6850 ;
      RECT 99.8350 240.1150 119.5000 240.6850 ;
      RECT 20.5000 240.1150 99.2650 240.6850 ;
      RECT 900.5000 238.8850 999.5000 240.1150 ;
      RECT 20.5000 238.8850 119.5000 240.1150 ;
      RECT 920.5700 238.3150 999.5000 238.8850 ;
      RECT 900.5000 238.3150 920.0000 238.8850 ;
      RECT 99.8350 238.3150 119.5000 238.8850 ;
      RECT 20.5000 238.3150 99.2650 238.8850 ;
      RECT 900.5000 237.0850 999.5000 238.3150 ;
      RECT 20.5000 237.0850 119.5000 238.3150 ;
      RECT 920.5700 236.5150 999.5000 237.0850 ;
      RECT 900.5000 236.5150 920.0000 237.0850 ;
      RECT 99.8350 236.5150 119.5000 237.0850 ;
      RECT 20.5000 236.5150 99.2650 237.0850 ;
      RECT 900.5000 235.2850 999.5000 236.5150 ;
      RECT 20.5000 235.2850 119.5000 236.5150 ;
      RECT 920.5700 234.7150 999.5000 235.2850 ;
      RECT 900.5000 234.7150 920.0000 235.2850 ;
      RECT 99.8350 234.7150 119.5000 235.2850 ;
      RECT 20.5000 234.7150 99.2650 235.2850 ;
      RECT 900.5000 233.4850 999.5000 234.7150 ;
      RECT 20.5000 233.4850 119.5000 234.7150 ;
      RECT 920.5700 232.9150 999.5000 233.4850 ;
      RECT 900.5000 232.9150 920.0000 233.4850 ;
      RECT 99.8350 232.9150 119.5000 233.4850 ;
      RECT 20.5000 232.9150 99.2650 233.4850 ;
      RECT 900.5000 231.6850 999.5000 232.9150 ;
      RECT 20.5000 231.6850 119.5000 232.9150 ;
      RECT 920.5700 231.1150 999.5000 231.6850 ;
      RECT 900.5000 231.1150 920.0000 231.6850 ;
      RECT 99.8350 231.1150 119.5000 231.6850 ;
      RECT 20.5000 231.1150 99.2650 231.6850 ;
      RECT 900.5000 229.8850 999.5000 231.1150 ;
      RECT 20.5000 229.8850 119.5000 231.1150 ;
      RECT 920.5700 229.3150 999.5000 229.8850 ;
      RECT 900.5000 229.3150 920.0000 229.8850 ;
      RECT 99.8350 229.3150 119.5000 229.8850 ;
      RECT 20.5000 229.3150 99.2650 229.8850 ;
      RECT 900.5000 228.0850 999.5000 229.3150 ;
      RECT 20.5000 228.0850 119.5000 229.3150 ;
      RECT 920.5700 227.5150 999.5000 228.0850 ;
      RECT 900.5000 227.5150 920.0000 228.0850 ;
      RECT 99.8350 227.5150 119.5000 228.0850 ;
      RECT 20.5000 227.5150 99.2650 228.0850 ;
      RECT 900.5000 226.2850 999.5000 227.5150 ;
      RECT 20.5000 226.2850 119.5000 227.5150 ;
      RECT 920.5700 225.7150 999.5000 226.2850 ;
      RECT 900.5000 225.7150 920.0000 226.2850 ;
      RECT 99.8350 225.7150 119.5000 226.2850 ;
      RECT 20.5000 225.7150 99.2650 226.2850 ;
      RECT 900.5000 224.4850 999.5000 225.7150 ;
      RECT 20.5000 224.4850 119.5000 225.7150 ;
      RECT 920.5700 223.9150 999.5000 224.4850 ;
      RECT 900.5000 223.9150 920.0000 224.4850 ;
      RECT 99.8350 223.9150 119.5000 224.4850 ;
      RECT 20.5000 223.9150 99.2650 224.4850 ;
      RECT 900.5000 222.6850 999.5000 223.9150 ;
      RECT 20.5000 222.6850 119.5000 223.9150 ;
      RECT 920.5700 222.1150 999.5000 222.6850 ;
      RECT 900.5000 222.1150 920.0000 222.6850 ;
      RECT 99.8350 222.1150 119.5000 222.6850 ;
      RECT 20.5000 222.1150 99.2650 222.6850 ;
      RECT 900.5000 220.8850 999.5000 222.1150 ;
      RECT 20.5000 220.8850 119.5000 222.1150 ;
      RECT 920.5700 220.3150 999.5000 220.8850 ;
      RECT 900.5000 220.3150 920.0000 220.8850 ;
      RECT 99.8350 220.3150 119.5000 220.8850 ;
      RECT 20.5000 220.3150 99.2650 220.8850 ;
      RECT 900.5000 219.0850 999.5000 220.3150 ;
      RECT 20.5000 219.0850 119.5000 220.3150 ;
      RECT 920.5700 218.5150 999.5000 219.0850 ;
      RECT 900.5000 218.5150 920.0000 219.0850 ;
      RECT 99.8350 218.5150 119.5000 219.0850 ;
      RECT 20.5000 218.5150 99.2650 219.0850 ;
      RECT 900.5000 217.2850 999.5000 218.5150 ;
      RECT 20.5000 217.2850 119.5000 218.5150 ;
      RECT 920.5700 216.7150 999.5000 217.2850 ;
      RECT 900.5000 216.7150 920.0000 217.2850 ;
      RECT 99.8350 216.7150 119.5000 217.2850 ;
      RECT 20.5000 216.7150 99.2650 217.2850 ;
      RECT 900.5000 215.4850 999.5000 216.7150 ;
      RECT 20.5000 215.4850 119.5000 216.7150 ;
      RECT 920.5700 214.9150 999.5000 215.4850 ;
      RECT 900.5000 214.9150 920.0000 215.4850 ;
      RECT 99.8350 214.9150 119.5000 215.4850 ;
      RECT 20.5000 214.9150 99.2650 215.4850 ;
      RECT 900.5000 213.6850 999.5000 214.9150 ;
      RECT 20.5000 213.6850 119.5000 214.9150 ;
      RECT 920.5700 213.1150 999.5000 213.6850 ;
      RECT 900.5000 213.1150 920.0000 213.6850 ;
      RECT 99.8350 213.1150 119.5000 213.6850 ;
      RECT 20.5000 213.1150 99.2650 213.6850 ;
      RECT 900.5000 211.8850 999.5000 213.1150 ;
      RECT 20.5000 211.8850 119.5000 213.1150 ;
      RECT 920.5700 211.3150 999.5000 211.8850 ;
      RECT 900.5000 211.3150 920.0000 211.8850 ;
      RECT 99.8350 211.3150 119.5000 211.8850 ;
      RECT 20.5000 211.3150 99.2650 211.8850 ;
      RECT 900.5000 210.0850 999.5000 211.3150 ;
      RECT 20.5000 210.0850 119.5000 211.3150 ;
      RECT 920.5700 209.5150 999.5000 210.0850 ;
      RECT 900.5000 209.5150 920.0000 210.0850 ;
      RECT 99.8350 209.5150 119.5000 210.0850 ;
      RECT 20.5000 209.5150 99.2650 210.0850 ;
      RECT 900.5000 208.2850 999.5000 209.5150 ;
      RECT 20.5000 208.2850 119.5000 209.5150 ;
      RECT 920.5700 207.7150 999.5000 208.2850 ;
      RECT 900.5000 207.7150 920.0000 208.2850 ;
      RECT 99.8350 207.7150 119.5000 208.2850 ;
      RECT 20.5000 207.7150 99.2650 208.2850 ;
      RECT 900.5000 206.4850 999.5000 207.7150 ;
      RECT 20.5000 206.4850 119.5000 207.7150 ;
      RECT 920.5700 205.9150 999.5000 206.4850 ;
      RECT 900.5000 205.9150 920.0000 206.4850 ;
      RECT 99.8350 205.9150 119.5000 206.4850 ;
      RECT 20.5000 205.9150 99.2650 206.4850 ;
      RECT 900.5000 204.6850 999.5000 205.9150 ;
      RECT 20.5000 204.6850 119.5000 205.9150 ;
      RECT 920.5700 204.1150 999.5000 204.6850 ;
      RECT 900.5000 204.1150 920.0000 204.6850 ;
      RECT 99.8350 204.1150 119.5000 204.6850 ;
      RECT 20.5000 204.1150 99.2650 204.6850 ;
      RECT 900.5000 202.8850 999.5000 204.1150 ;
      RECT 20.5000 202.8850 119.5000 204.1150 ;
      RECT 920.5700 202.3150 999.5000 202.8850 ;
      RECT 900.5000 202.3150 920.0000 202.8850 ;
      RECT 99.8350 202.3150 119.5000 202.8850 ;
      RECT 20.5000 202.3150 99.2650 202.8850 ;
      RECT 900.5000 201.0850 999.5000 202.3150 ;
      RECT 20.5000 201.0850 119.5000 202.3150 ;
      RECT 920.5700 200.5150 999.5000 201.0850 ;
      RECT 900.5000 200.5150 920.0000 201.0850 ;
      RECT 99.8350 200.5150 119.5000 201.0850 ;
      RECT 20.5000 200.5150 99.2650 201.0850 ;
      RECT 900.5000 199.2850 999.5000 200.5150 ;
      RECT 20.5000 199.2850 119.5000 200.5150 ;
      RECT 920.5700 198.7150 999.5000 199.2850 ;
      RECT 900.5000 198.7150 920.0000 199.2850 ;
      RECT 99.8350 198.7150 119.5000 199.2850 ;
      RECT 20.5000 198.7150 99.2650 199.2850 ;
      RECT 900.5000 197.4850 999.5000 198.7150 ;
      RECT 20.5000 197.4850 119.5000 198.7150 ;
      RECT 920.5700 196.9150 999.5000 197.4850 ;
      RECT 900.5000 196.9150 920.0000 197.4850 ;
      RECT 99.8350 196.9150 119.5000 197.4850 ;
      RECT 20.5000 196.9150 99.2650 197.4850 ;
      RECT 900.5000 195.6850 999.5000 196.9150 ;
      RECT 20.5000 195.6850 119.5000 196.9150 ;
      RECT 920.5700 195.1150 999.5000 195.6850 ;
      RECT 900.5000 195.1150 920.0000 195.6850 ;
      RECT 99.8350 195.1150 119.5000 195.6850 ;
      RECT 20.5000 195.1150 99.2650 195.6850 ;
      RECT 900.5000 193.8850 999.5000 195.1150 ;
      RECT 20.5000 193.8850 119.5000 195.1150 ;
      RECT 920.5700 193.3150 999.5000 193.8850 ;
      RECT 900.5000 193.3150 920.0000 193.8850 ;
      RECT 99.8350 193.3150 119.5000 193.8850 ;
      RECT 20.5000 193.3150 99.2650 193.8850 ;
      RECT 900.5000 192.0850 999.5000 193.3150 ;
      RECT 20.5000 192.0850 119.5000 193.3150 ;
      RECT 920.5700 191.5150 999.5000 192.0850 ;
      RECT 900.5000 191.5150 920.0000 192.0850 ;
      RECT 99.8350 191.5150 119.5000 192.0850 ;
      RECT 20.5000 191.5150 99.2650 192.0850 ;
      RECT 900.5000 190.2850 999.5000 191.5150 ;
      RECT 20.5000 190.2850 119.5000 191.5150 ;
      RECT 920.5700 189.7150 999.5000 190.2850 ;
      RECT 900.5000 189.7150 920.0000 190.2850 ;
      RECT 99.8350 189.7150 119.5000 190.2850 ;
      RECT 20.5000 189.7150 99.2650 190.2850 ;
      RECT 900.5000 188.4850 999.5000 189.7150 ;
      RECT 20.5000 188.4850 119.5000 189.7150 ;
      RECT 920.5700 187.9150 999.5000 188.4850 ;
      RECT 900.5000 187.9150 920.0000 188.4850 ;
      RECT 99.8350 187.9150 119.5000 188.4850 ;
      RECT 20.5000 187.9150 99.2650 188.4850 ;
      RECT 900.5000 186.6850 999.5000 187.9150 ;
      RECT 20.5000 186.6850 119.5000 187.9150 ;
      RECT 920.5700 186.1150 999.5000 186.6850 ;
      RECT 900.5000 186.1150 920.0000 186.6850 ;
      RECT 99.8350 186.1150 119.5000 186.6850 ;
      RECT 20.5000 186.1150 99.2650 186.6850 ;
      RECT 900.5000 184.8850 999.5000 186.1150 ;
      RECT 20.5000 184.8850 119.5000 186.1150 ;
      RECT 920.5700 184.3150 999.5000 184.8850 ;
      RECT 900.5000 184.3150 920.0000 184.8850 ;
      RECT 99.8350 184.3150 119.5000 184.8850 ;
      RECT 20.5000 184.3150 99.2650 184.8850 ;
      RECT 900.5000 183.0850 999.5000 184.3150 ;
      RECT 20.5000 183.0850 119.5000 184.3150 ;
      RECT 920.5700 182.5150 999.5000 183.0850 ;
      RECT 900.5000 182.5150 920.0000 183.0850 ;
      RECT 99.8350 182.5150 119.5000 183.0850 ;
      RECT 20.5000 182.5150 99.2650 183.0850 ;
      RECT 900.5000 181.2850 999.5000 182.5150 ;
      RECT 20.5000 181.2850 119.5000 182.5150 ;
      RECT 920.5700 180.7150 999.5000 181.2850 ;
      RECT 900.5000 180.7150 920.0000 181.2850 ;
      RECT 99.8350 180.7150 119.5000 181.2850 ;
      RECT 20.5000 180.7150 99.2650 181.2850 ;
      RECT 900.5000 179.4850 999.5000 180.7150 ;
      RECT 20.5000 179.4850 119.5000 180.7150 ;
      RECT 920.5700 178.9150 999.5000 179.4850 ;
      RECT 900.5000 178.9150 920.0000 179.4850 ;
      RECT 99.8350 178.9150 119.5000 179.4850 ;
      RECT 20.5000 178.9150 99.2650 179.4850 ;
      RECT 900.5000 177.6850 999.5000 178.9150 ;
      RECT 20.5000 177.6850 119.5000 178.9150 ;
      RECT 920.5700 177.1150 999.5000 177.6850 ;
      RECT 900.5000 177.1150 920.0000 177.6850 ;
      RECT 99.8350 177.1150 119.5000 177.6850 ;
      RECT 20.5000 177.1150 99.2650 177.6850 ;
      RECT 900.5000 175.8850 999.5000 177.1150 ;
      RECT 20.5000 175.8850 119.5000 177.1150 ;
      RECT 920.5700 175.3150 999.5000 175.8850 ;
      RECT 900.5000 175.3150 920.0000 175.8850 ;
      RECT 99.8350 175.3150 119.5000 175.8850 ;
      RECT 20.5000 175.3150 99.2650 175.8850 ;
      RECT 900.5000 174.0850 999.5000 175.3150 ;
      RECT 20.5000 174.0850 119.5000 175.3150 ;
      RECT 920.5700 173.5150 999.5000 174.0850 ;
      RECT 900.5000 173.5150 920.0000 174.0850 ;
      RECT 99.8350 173.5150 119.5000 174.0850 ;
      RECT 20.5000 173.5150 99.2650 174.0850 ;
      RECT 900.5000 172.2850 999.5000 173.5150 ;
      RECT 20.5000 172.2850 119.5000 173.5150 ;
      RECT 920.5700 171.7150 999.5000 172.2850 ;
      RECT 900.5000 171.7150 920.0000 172.2850 ;
      RECT 99.8350 171.7150 119.5000 172.2850 ;
      RECT 20.5000 171.7150 99.2650 172.2850 ;
      RECT 900.5000 170.4850 999.5000 171.7150 ;
      RECT 20.5000 170.4850 119.5000 171.7150 ;
      RECT 920.5700 169.9150 999.5000 170.4850 ;
      RECT 900.5000 169.9150 920.0000 170.4850 ;
      RECT 99.8350 169.9150 119.5000 170.4850 ;
      RECT 20.5000 169.9150 99.2650 170.4850 ;
      RECT 900.5000 168.6850 999.5000 169.9150 ;
      RECT 20.5000 168.6850 119.5000 169.9150 ;
      RECT 920.5700 168.1150 999.5000 168.6850 ;
      RECT 900.5000 168.1150 920.0000 168.6850 ;
      RECT 99.8350 168.1150 119.5000 168.6850 ;
      RECT 20.5000 168.1150 99.2650 168.6850 ;
      RECT 900.5000 166.8850 999.5000 168.1150 ;
      RECT 20.5000 166.8850 119.5000 168.1150 ;
      RECT 920.5700 166.3150 999.5000 166.8850 ;
      RECT 900.5000 166.3150 920.0000 166.8850 ;
      RECT 99.8350 166.3150 119.5000 166.8850 ;
      RECT 20.5000 166.3150 99.2650 166.8850 ;
      RECT 900.5000 165.0850 999.5000 166.3150 ;
      RECT 20.5000 165.0850 119.5000 166.3150 ;
      RECT 920.5700 164.5150 999.5000 165.0850 ;
      RECT 900.5000 164.5150 920.0000 165.0850 ;
      RECT 99.8350 164.5150 119.5000 165.0850 ;
      RECT 20.5000 164.5150 99.2650 165.0850 ;
      RECT 900.5000 163.2850 999.5000 164.5150 ;
      RECT 20.5000 163.2850 119.5000 164.5150 ;
      RECT 920.5700 162.7150 999.5000 163.2850 ;
      RECT 900.5000 162.7150 920.0000 163.2850 ;
      RECT 99.8350 162.7150 119.5000 163.2850 ;
      RECT 20.5000 162.7150 99.2650 163.2850 ;
      RECT 900.5000 161.4850 999.5000 162.7150 ;
      RECT 20.5000 161.4850 119.5000 162.7150 ;
      RECT 920.5700 160.9150 999.5000 161.4850 ;
      RECT 900.5000 160.9150 920.0000 161.4850 ;
      RECT 99.8350 160.9150 119.5000 161.4850 ;
      RECT 20.5000 160.9150 99.2650 161.4850 ;
      RECT 900.5000 159.6850 999.5000 160.9150 ;
      RECT 20.5000 159.6850 119.5000 160.9150 ;
      RECT 920.5700 159.1150 999.5000 159.6850 ;
      RECT 900.5000 159.1150 920.0000 159.6850 ;
      RECT 99.8350 159.1150 119.5000 159.6850 ;
      RECT 20.5000 159.1150 99.2650 159.6850 ;
      RECT 900.5000 157.8850 999.5000 159.1150 ;
      RECT 20.5000 157.8850 119.5000 159.1150 ;
      RECT 920.5700 157.3150 999.5000 157.8850 ;
      RECT 900.5000 157.3150 920.0000 157.8850 ;
      RECT 99.8350 157.3150 119.5000 157.8850 ;
      RECT 20.5000 157.3150 99.2650 157.8850 ;
      RECT 900.5000 156.0850 999.5000 157.3150 ;
      RECT 20.5000 156.0850 119.5000 157.3150 ;
      RECT 920.5700 155.5150 999.5000 156.0850 ;
      RECT 900.5000 155.5150 920.0000 156.0850 ;
      RECT 99.8350 155.5150 119.5000 156.0850 ;
      RECT 20.5000 155.5150 99.2650 156.0850 ;
      RECT 900.5000 154.2850 999.5000 155.5150 ;
      RECT 20.5000 154.2850 119.5000 155.5150 ;
      RECT 920.5700 153.7150 999.5000 154.2850 ;
      RECT 900.5000 153.7150 920.0000 154.2850 ;
      RECT 99.8350 153.7150 119.5000 154.2850 ;
      RECT 20.5000 153.7150 99.2650 154.2850 ;
      RECT 900.5000 152.4850 999.5000 153.7150 ;
      RECT 20.5000 152.4850 119.5000 153.7150 ;
      RECT 920.5700 151.9150 999.5000 152.4850 ;
      RECT 900.5000 151.9150 920.0000 152.4850 ;
      RECT 99.8350 151.9150 119.5000 152.4850 ;
      RECT 20.5000 151.9150 99.2650 152.4850 ;
      RECT 900.5000 150.6850 999.5000 151.9150 ;
      RECT 20.5000 150.6850 119.5000 151.9150 ;
      RECT 920.5700 150.1150 999.5000 150.6850 ;
      RECT 900.5000 150.1150 920.0000 150.6850 ;
      RECT 99.8350 150.1150 119.5000 150.6850 ;
      RECT 20.5000 150.1150 99.2650 150.6850 ;
      RECT 900.5000 148.8850 999.5000 150.1150 ;
      RECT 20.5000 148.8850 119.5000 150.1150 ;
      RECT 920.5700 148.3150 999.5000 148.8850 ;
      RECT 900.5000 148.3150 920.0000 148.8850 ;
      RECT 99.8350 148.3150 119.5000 148.8850 ;
      RECT 20.5000 148.3150 99.2650 148.8850 ;
      RECT 900.5000 147.0850 999.5000 148.3150 ;
      RECT 20.5000 147.0850 119.5000 148.3150 ;
      RECT 920.5700 146.5150 999.5000 147.0850 ;
      RECT 900.5000 146.5150 920.0000 147.0850 ;
      RECT 99.8350 146.5150 119.5000 147.0850 ;
      RECT 20.5000 146.5150 99.2650 147.0850 ;
      RECT 900.5000 145.2850 999.5000 146.5150 ;
      RECT 20.5000 145.2850 119.5000 146.5150 ;
      RECT 920.5700 144.7150 999.5000 145.2850 ;
      RECT 900.5000 144.7150 920.0000 145.2850 ;
      RECT 99.8350 144.7150 119.5000 145.2850 ;
      RECT 20.5000 144.7150 99.2650 145.2850 ;
      RECT 900.5000 143.4850 999.5000 144.7150 ;
      RECT 20.5000 143.4850 119.5000 144.7150 ;
      RECT 920.5700 142.9150 999.5000 143.4850 ;
      RECT 900.5000 142.9150 920.0000 143.4850 ;
      RECT 99.8350 142.9150 119.5000 143.4850 ;
      RECT 20.5000 142.9150 99.2650 143.4850 ;
      RECT 900.5000 141.6850 999.5000 142.9150 ;
      RECT 20.5000 141.6850 119.5000 142.9150 ;
      RECT 920.5700 141.1150 999.5000 141.6850 ;
      RECT 900.5000 141.1150 920.0000 141.6850 ;
      RECT 99.8350 141.1150 119.5000 141.6850 ;
      RECT 20.5000 141.1150 99.2650 141.6850 ;
      RECT 900.5000 139.8850 999.5000 141.1150 ;
      RECT 20.5000 139.8850 119.5000 141.1150 ;
      RECT 920.5700 139.3150 999.5000 139.8850 ;
      RECT 900.5000 139.3150 920.0000 139.8850 ;
      RECT 99.8350 139.3150 119.5000 139.8850 ;
      RECT 20.5000 139.3150 99.2650 139.8850 ;
      RECT 900.5000 138.0850 999.5000 139.3150 ;
      RECT 20.5000 138.0850 119.5000 139.3150 ;
      RECT 920.5700 137.5150 999.5000 138.0850 ;
      RECT 900.5000 137.5150 920.0000 138.0850 ;
      RECT 99.8350 137.5150 119.5000 138.0850 ;
      RECT 20.5000 137.5150 99.2650 138.0850 ;
      RECT 900.5000 136.2850 999.5000 137.5150 ;
      RECT 20.5000 136.2850 119.5000 137.5150 ;
      RECT 920.5700 135.7150 999.5000 136.2850 ;
      RECT 900.5000 135.7150 920.0000 136.2850 ;
      RECT 99.8350 135.7150 119.5000 136.2850 ;
      RECT 20.5000 135.7150 99.2650 136.2850 ;
      RECT 900.5000 134.4850 999.5000 135.7150 ;
      RECT 20.5000 134.4850 119.5000 135.7150 ;
      RECT 920.5700 133.9150 999.5000 134.4850 ;
      RECT 900.5000 133.9150 920.0000 134.4850 ;
      RECT 99.8350 133.9150 119.5000 134.4850 ;
      RECT 20.5000 133.9150 99.2650 134.4850 ;
      RECT 900.5000 132.6850 999.5000 133.9150 ;
      RECT 20.5000 132.6850 119.5000 133.9150 ;
      RECT 920.5700 132.1150 999.5000 132.6850 ;
      RECT 900.5000 132.1150 920.0000 132.6850 ;
      RECT 99.8350 132.1150 119.5000 132.6850 ;
      RECT 20.5000 132.1150 99.2650 132.6850 ;
      RECT 900.5000 130.8850 999.5000 132.1150 ;
      RECT 20.5000 130.8850 119.5000 132.1150 ;
      RECT 920.5700 130.3150 999.5000 130.8850 ;
      RECT 900.5000 130.3150 920.0000 130.8850 ;
      RECT 99.8350 130.3150 119.5000 130.8850 ;
      RECT 20.5000 130.3150 99.2650 130.8850 ;
      RECT 900.5000 129.0850 999.5000 130.3150 ;
      RECT 20.5000 129.0850 119.5000 130.3150 ;
      RECT 920.5700 128.5150 999.5000 129.0850 ;
      RECT 900.5000 128.5150 920.0000 129.0850 ;
      RECT 99.8350 128.5150 119.5000 129.0850 ;
      RECT 20.5000 128.5150 99.2650 129.0850 ;
      RECT 900.5000 127.2850 999.5000 128.5150 ;
      RECT 20.5000 127.2850 119.5000 128.5150 ;
      RECT 920.5700 126.7150 999.5000 127.2850 ;
      RECT 900.5000 126.7150 920.0000 127.2850 ;
      RECT 99.8350 126.7150 119.5000 127.2850 ;
      RECT 20.5000 126.7150 99.2650 127.2850 ;
      RECT 900.5000 125.4850 999.5000 126.7150 ;
      RECT 20.5000 125.4850 119.5000 126.7150 ;
      RECT 920.5700 124.9150 999.5000 125.4850 ;
      RECT 900.5000 124.9150 920.0000 125.4850 ;
      RECT 99.8350 124.9150 119.5000 125.4850 ;
      RECT 20.5000 124.9150 99.2650 125.4850 ;
      RECT 900.5000 123.6850 999.5000 124.9150 ;
      RECT 20.5000 123.6850 119.5000 124.9150 ;
      RECT 920.5700 123.1150 999.5000 123.6850 ;
      RECT 900.5000 123.1150 920.0000 123.6850 ;
      RECT 99.8350 123.1150 119.5000 123.6850 ;
      RECT 20.5000 123.1150 99.2650 123.6850 ;
      RECT 900.5000 121.8850 999.5000 123.1150 ;
      RECT 20.5000 121.8850 119.5000 123.1150 ;
      RECT 920.5700 121.3150 999.5000 121.8850 ;
      RECT 900.5000 121.3150 920.0000 121.8850 ;
      RECT 99.8350 121.3150 119.5000 121.8850 ;
      RECT 20.5000 121.3150 99.2650 121.8850 ;
      RECT 900.5000 120.0850 999.5000 121.3150 ;
      RECT 20.5000 120.0850 119.5000 121.3150 ;
      RECT 920.5700 119.5150 999.5000 120.0850 ;
      RECT 900.5000 119.5150 920.0000 120.0850 ;
      RECT 99.8350 119.5150 119.5000 120.0850 ;
      RECT 20.5000 119.5150 99.2650 120.0850 ;
      RECT 900.5000 118.2850 999.5000 119.5150 ;
      RECT 20.5000 118.2850 119.5000 119.5150 ;
      RECT 920.5700 117.7150 999.5000 118.2850 ;
      RECT 900.5000 117.7150 920.0000 118.2850 ;
      RECT 99.8350 117.7150 119.5000 118.2850 ;
      RECT 20.5000 117.7150 99.2650 118.2850 ;
      RECT 900.5000 116.4850 999.5000 117.7150 ;
      RECT 20.5000 116.4850 119.5000 117.7150 ;
      RECT 920.5700 115.9150 999.5000 116.4850 ;
      RECT 900.5000 115.9150 920.0000 116.4850 ;
      RECT 99.8350 115.9150 119.5000 116.4850 ;
      RECT 20.5000 115.9150 99.2650 116.4850 ;
      RECT 900.5000 114.6850 999.5000 115.9150 ;
      RECT 20.5000 114.6850 119.5000 115.9150 ;
      RECT 920.5700 114.1150 999.5000 114.6850 ;
      RECT 900.5000 114.1150 920.0000 114.6850 ;
      RECT 99.8350 114.1150 119.5000 114.6850 ;
      RECT 20.5000 114.1150 99.2650 114.6850 ;
      RECT 900.5000 112.8850 999.5000 114.1150 ;
      RECT 20.5000 112.8850 119.5000 114.1150 ;
      RECT 920.5700 112.3150 999.5000 112.8850 ;
      RECT 900.5000 112.3150 920.0000 112.8850 ;
      RECT 99.8350 112.3150 119.5000 112.8850 ;
      RECT 20.5000 112.3150 99.2650 112.8850 ;
      RECT 900.5000 111.0850 999.5000 112.3150 ;
      RECT 20.5000 111.0850 119.5000 112.3150 ;
      RECT 920.5700 110.5150 999.5000 111.0850 ;
      RECT 900.5000 110.5150 920.0000 111.0850 ;
      RECT 99.8350 110.5150 119.5000 111.0850 ;
      RECT 20.5000 110.5150 99.2650 111.0850 ;
      RECT 900.5000 109.2850 999.5000 110.5150 ;
      RECT 20.5000 109.2850 119.5000 110.5150 ;
      RECT 920.5700 108.7150 999.5000 109.2850 ;
      RECT 900.5000 108.7150 920.0000 109.2850 ;
      RECT 99.8350 108.7150 119.5000 109.2850 ;
      RECT 20.5000 108.7150 99.2650 109.2850 ;
      RECT 900.5000 107.4850 999.5000 108.7150 ;
      RECT 20.5000 107.4850 119.5000 108.7150 ;
      RECT 920.5700 106.9150 999.5000 107.4850 ;
      RECT 900.5000 106.9150 920.0000 107.4850 ;
      RECT 99.8350 106.9150 119.5000 107.4850 ;
      RECT 20.5000 106.9150 99.2650 107.4850 ;
      RECT 900.5000 105.6850 999.5000 106.9150 ;
      RECT 20.5000 105.6850 119.5000 106.9150 ;
      RECT 920.5700 105.1150 999.5000 105.6850 ;
      RECT 900.5000 105.1150 920.0000 105.6850 ;
      RECT 99.8350 105.1150 119.5000 105.6850 ;
      RECT 20.5000 105.1150 99.2650 105.6850 ;
      RECT 900.5000 103.8850 999.5000 105.1150 ;
      RECT 20.5000 103.8850 119.5000 105.1150 ;
      RECT 920.5700 103.3150 999.5000 103.8850 ;
      RECT 900.5000 103.3150 920.0000 103.8850 ;
      RECT 99.8350 103.3150 119.5000 103.8850 ;
      RECT 20.5000 103.3150 99.2650 103.8850 ;
      RECT 900.5000 102.0850 999.5000 103.3150 ;
      RECT 20.5000 102.0850 119.5000 103.3150 ;
      RECT 920.5700 101.5150 999.5000 102.0850 ;
      RECT 900.5000 101.5150 920.0000 102.0850 ;
      RECT 99.8350 101.5150 119.5000 102.0850 ;
      RECT 20.5000 101.5150 99.2650 102.0850 ;
      RECT 900.5000 100.2850 999.5000 101.5150 ;
      RECT 20.5000 100.2850 119.5000 101.5150 ;
      RECT 920.5700 99.7150 999.5000 100.2850 ;
      RECT 900.5000 99.7150 920.0000 100.2850 ;
      RECT 99.8350 99.7150 119.5000 100.2850 ;
      RECT 20.5000 99.7150 99.2650 100.2850 ;
      RECT 1002.5000 9.5000 1007.5000 1610.5000 ;
      RECT 900.5000 9.5000 999.5000 99.7150 ;
      RECT 892.5000 9.5000 897.5000 1610.5000 ;
      RECT 790.5000 9.5000 889.5000 1610.5000 ;
      RECT 782.5000 9.5000 787.5000 1610.5000 ;
      RECT 680.5000 9.5000 779.5000 1610.5000 ;
      RECT 672.5000 9.5000 677.5000 1610.5000 ;
      RECT 570.5000 9.5000 669.5000 1610.5000 ;
      RECT 562.5000 9.5000 567.5000 1610.5000 ;
      RECT 460.5000 9.5000 559.5000 1610.5000 ;
      RECT 452.5000 9.5000 457.5000 1610.5000 ;
      RECT 350.5000 9.5000 449.5000 1610.5000 ;
      RECT 342.5000 9.5000 347.5000 1610.5000 ;
      RECT 240.5000 9.5000 339.5000 1610.5000 ;
      RECT 232.5000 9.5000 237.5000 1610.5000 ;
      RECT 130.5000 9.5000 229.5000 1610.5000 ;
      RECT 122.5000 9.5000 127.5000 1610.5000 ;
      RECT 20.5000 9.5000 119.5000 99.7150 ;
      RECT 12.5000 9.5000 17.5000 1610.5000 ;
      RECT 0.0000 9.5000 9.5000 1610.5000 ;
      RECT 1010.5000 9.3350 1020.0000 1610.5000 ;
      RECT 900.5000 9.3350 1007.5000 9.5000 ;
      RECT 790.5000 9.3350 897.5000 9.5000 ;
      RECT 680.5000 9.3350 787.5000 9.5000 ;
      RECT 570.5000 9.3350 677.5000 9.5000 ;
      RECT 460.5000 9.3350 567.5000 9.5000 ;
      RECT 350.5000 9.3350 457.5000 9.5000 ;
      RECT 240.5000 9.3350 347.5000 9.5000 ;
      RECT 130.5000 9.3350 237.5000 9.5000 ;
      RECT 20.5000 9.3350 127.5000 9.5000 ;
      RECT 0.0000 9.3350 17.5000 9.5000 ;
      RECT 0.0000 0.0000 1020.0000 9.3350 ;
  END
END core

END LIBRARY
